* PEX netlist file	Mon May  2 16:35:55 2022	and_2
* icv_netlist Version RHEL64 S-2021.06-SP2.6831572 2021/08/30
*.UNIT=4000

* Hierarchy Level 0

* Top of hierarchy  cell=and_2
.subckt and_2 A 3 Z GND! VDD! B 8
*.floating_nets _GENERATED_9 _GENERATED_10 _GENERATED_11 _GENERATED_12
MM1 Z 3 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2450 $Y=1254  $PIN_XY=2480,1082,2450,1254,2420,1082 $DEVICE_ID=1001
MM2 3 A 8 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=1946 $Y=972  $PIN_XY=(1976,1082,1976,912),1946,972,(1916,1082,1916,912) $DEVICE_ID=1001
MM3 8 B GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=1778 $Y=1167  $PIN_XY=(1808,1082,1808,912),1778,1167,(1748,1082,1748,912) $DEVICE_ID=1001
MM4 Z 3 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2450 $Y=1254  $PIN_XY=(2480,1422,2480,1252),2450,1254,(2420,1422,2420,1252) $DEVICE_ID=1003
MM5 3 A VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2114 $Y=1355  $PIN_XY=(2144,1422,2144,1252),2114,1355,(2084,1422,2084,1252) $DEVICE_ID=1003
MM6 3 B VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1778 $Y=1167  $PIN_XY=(1808,1422,1808,1252),1778,1167,(1748,1422,1748,1252) $DEVICE_ID=1003
.ends and_2
