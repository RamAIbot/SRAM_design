* PEX netlist file	Wed Apr 20 01:54:39 2022	rowdecoder
* icv_netlist Version RHEL64 S-2021.06-SP2.6831572 2021/08/30
*.UNIT=4000

* Hierarchy Level 1
.subckt inv_2 2 3 4 5 6 7
*.floating_nets _GENERATED_8
MM1 3 2 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=0 $Y=170  $PIN_XY=30,0,0,170,-30,0 $DEVICE_ID=1001
MM2 3 2 5 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=0 $Y=170  $PIN_XY=(30,340,30,170),0,170,(-30,340,-30,170) $DEVICE_ID=1003
.ends inv_2
.subckt nor_5 2 3 4 5 6 7 8 9 10 11
*.floating_nets _GENERATED_12 _GENERATED_13
.ends nor_5

* Hierarchy Level 0

* Top of hierarchy  cell=rowdecoder
.subckt rowdecoder A<4> A<3> A<2> 5 6 7 WL<0> WL<1> WL<2> WL<3> WL<4>
+	WL<5> WL<6> WL<7> VDD! GND!
*.floating_nets 8 9 _GENERATED_153 _GENERATED_154 _GENERATED_155 _GENERATED_156 _GENERATED_157 _GENERATED_158 _GENERATED_159 _GENERATED_160 _GENERATED_161
*+	_GENERATED_162 _GENERATED_163 _GENERATED_164
MM1 WL<0> A<3> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3722 $Y=9152  $PIN_XY=3752,9152,3722,9152,3692,9152 $DEVICE_ID=1001
MM2 WL<1> A<3> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3722 $Y=8004  $PIN_XY=3752,8004,3722,8004,3692,8004 $DEVICE_ID=1001
MM3 WL<2> 6 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3722 $Y=6854  $PIN_XY=3752,6854,3722,6854,3692,6854 $DEVICE_ID=1001
MM4 WL<3> 6 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3722 $Y=5706  $PIN_XY=3752,5706,3722,5706,3692,5706 $DEVICE_ID=1001
MM5 WL<4> A<3> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3722 $Y=4558  $PIN_XY=3752,4558,3722,4558,3692,4558 $DEVICE_ID=1001
MM6 WL<5> A<3> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3722 $Y=3410  $PIN_XY=3752,3410,3722,3410,3692,3410 $DEVICE_ID=1001
MM7 WL<6> 6 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3722 $Y=2262  $PIN_XY=3752,2262,3722,2262,3692,2262 $DEVICE_ID=1001
MM8 WL<7> 6 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3722 $Y=1114  $PIN_XY=3752,1114,3722,1114,3692,1114 $DEVICE_ID=1001
MM9 WL<0> A<2> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3386 $Y=9350  $PIN_XY=3416,9152,3386,9350,3356,9152 $DEVICE_ID=1001
MM10 WL<1> 5 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3386 $Y=8202  $PIN_XY=3416,8004,3386,8202,3356,8004 $DEVICE_ID=1001
MM11 WL<2> A<2> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3386 $Y=7052  $PIN_XY=3416,6854,3386,7052,3356,6854 $DEVICE_ID=1001
MM12 WL<3> 5 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3386 $Y=5904  $PIN_XY=3416,5706,3386,5904,3356,5706 $DEVICE_ID=1001
MM13 WL<4> A<2> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3386 $Y=4756  $PIN_XY=3416,4558,3386,4756,3356,4558 $DEVICE_ID=1001
MM14 WL<5> 5 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3386 $Y=3608  $PIN_XY=3416,3410,3386,3608,3356,3410 $DEVICE_ID=1001
MM15 WL<6> A<2> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3386 $Y=2460  $PIN_XY=3416,2262,3386,2460,3356,2262 $DEVICE_ID=1001
MM16 WL<7> 5 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3386 $Y=1312  $PIN_XY=3416,1114,3386,1312,3356,1114 $DEVICE_ID=1001
MM17 WL<0> A<4> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3050 $Y=9350  $PIN_XY=3080,9152,3050,9350,3020,9152 $DEVICE_ID=1001
MM18 WL<1> A<4> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3050 $Y=8202  $PIN_XY=3080,8004,3050,8202,3020,8004 $DEVICE_ID=1001
MM19 WL<2> A<4> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3050 $Y=7052  $PIN_XY=3080,6854,3050,7052,3020,6854 $DEVICE_ID=1001
MM20 WL<3> A<4> GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3050 $Y=5904  $PIN_XY=3080,5706,3050,5904,3020,5706 $DEVICE_ID=1001
MM21 WL<4> 7 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3050 $Y=4756  $PIN_XY=3080,4558,3050,4756,3020,4558 $DEVICE_ID=1001
MM22 WL<5> 7 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3050 $Y=3608  $PIN_XY=3080,3410,3050,3608,3020,3410 $DEVICE_ID=1001
MM23 WL<6> 7 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3050 $Y=2460  $PIN_XY=3080,2262,3050,2460,3020,2262 $DEVICE_ID=1001
MM24 WL<7> 7 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3050 $Y=1312  $PIN_XY=3080,1114,3050,1312,3020,1114 $DEVICE_ID=1001
MM25 WL<0> A<2> 29 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3386 $Y=9350  $PIN_XY=(3416,9548,3416,9378),3386,9350,(3356,9548,3356,9378) $DEVICE_ID=1003
MM26 WL<1> 5 31 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3386 $Y=8202  $PIN_XY=(3416,8400,3416,8230),3386,8202,(3356,8400,3356,8230) $DEVICE_ID=1003
MM27 WL<2> A<2> 33 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3386 $Y=7052  $PIN_XY=(3416,7250,3416,7080),3386,7052,(3356,7250,3356,7080) $DEVICE_ID=1003
MM28 WL<3> 5 35 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3386 $Y=5904  $PIN_XY=(3416,6102,3416,5932),3386,5904,(3356,6102,3356,5932) $DEVICE_ID=1003
MM29 WL<4> A<2> 37 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3386 $Y=4756  $PIN_XY=(3416,4954,3416,4784),3386,4756,(3356,4954,3356,4784) $DEVICE_ID=1003
MM30 WL<5> 5 39 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3386 $Y=3608  $PIN_XY=(3416,3806,3416,3636),3386,3608,(3356,3806,3356,3636) $DEVICE_ID=1003
MM31 WL<6> A<2> 41 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3386 $Y=2460  $PIN_XY=(3416,2658,3416,2488),3386,2460,(3356,2658,3356,2488) $DEVICE_ID=1003
MM32 WL<7> 5 43 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3386 $Y=1312  $PIN_XY=(3416,1510,3416,1340),3386,1312,(3356,1510,3356,1340) $DEVICE_ID=1003
MM33 29 A<3> 28 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=3218 $Y=9450  $PIN_XY=(3248,9548,3248,9378),3218,9450,(3188,9548,3188,9378) $DEVICE_ID=1003
MM34 31 A<3> 30 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=3218 $Y=8302  $PIN_XY=(3248,8400,3248,8230),3218,8302,(3188,8400,3188,8230) $DEVICE_ID=1003
MM35 33 6 32 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=3218 $Y=7152  $PIN_XY=(3248,7250,3248,7080),3218,7152,(3188,7250,3188,7080) $DEVICE_ID=1003
MM36 35 6 34 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=3218 $Y=6004  $PIN_XY=(3248,6102,3248,5932),3218,6004,(3188,6102,3188,5932) $DEVICE_ID=1003
MM37 37 A<3> 36 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=3218 $Y=4856  $PIN_XY=(3248,4954,3248,4784),3218,4856,(3188,4954,3188,4784) $DEVICE_ID=1003
MM38 39 A<3> 38 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=3218 $Y=3708  $PIN_XY=(3248,3806,3248,3636),3218,3708,(3188,3806,3188,3636) $DEVICE_ID=1003
MM39 41 6 40 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=3218 $Y=2560  $PIN_XY=(3248,2658,3248,2488),3218,2560,(3188,2658,3188,2488) $DEVICE_ID=1003
MM40 43 6 42 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=3218 $Y=1412  $PIN_XY=(3248,1510,3248,1340),3218,1412,(3188,1510,3188,1340) $DEVICE_ID=1003
MM41 28 A<4> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3050 $Y=9350  $PIN_XY=(3080,9548,3080,9378),3050,9350,(3020,9548,3020,9378) $DEVICE_ID=1003
MM42 30 A<4> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3050 $Y=8202  $PIN_XY=(3080,8400,3080,8230),3050,8202,(3020,8400,3020,8230) $DEVICE_ID=1003
MM43 32 A<4> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3050 $Y=7052  $PIN_XY=(3080,7250,3080,7080),3050,7052,(3020,7250,3020,7080) $DEVICE_ID=1003
MM44 34 A<4> VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3050 $Y=5904  $PIN_XY=(3080,6102,3080,5932),3050,5904,(3020,6102,3020,5932) $DEVICE_ID=1003
MM45 36 7 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3050 $Y=4756  $PIN_XY=(3080,4954,3080,4784),3050,4756,(3020,4954,3020,4784) $DEVICE_ID=1003
MM46 38 7 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3050 $Y=3608  $PIN_XY=(3080,3806,3080,3636),3050,3608,(3020,3806,3020,3636) $DEVICE_ID=1003
MM47 40 7 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3050 $Y=2460  $PIN_XY=(3080,2658,3080,2488),3050,2460,(3020,2658,3020,2488) $DEVICE_ID=1003
MM48 42 7 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3050 $Y=1312  $PIN_XY=(3080,1510,3080,1340),3050,1312,(3020,1510,3020,1340) $DEVICE_ID=1003
XXFC9F1AD01 A<4> A<3> A<2> WL<0> GND! VDD! 28 29 20 VDD! nor_5 $T=3238 9162 0 0 $X=2824 $Y=8944
XXFC9F1AD02 A<4> A<3> 5 WL<1> GND! VDD! 30 31 21 VDD! nor_5 $T=3238 8014 0 0 $X=2824 $Y=7795
XXFC9F1AD03 A<4> 6 A<2> WL<2> GND! VDD! 32 33 22 VDD! nor_5 $T=3238 6864 0 0 $X=2824 $Y=6646
XXFC9F1AD04 A<4> 6 5 WL<3> GND! VDD! 34 35 23 VDD! nor_5 $T=3238 5716 0 0 $X=2824 $Y=5498
XXFC9F1AD05 7 A<3> A<2> WL<4> GND! VDD! 36 37 24 VDD! nor_5 $T=3238 4568 0 0 $X=2824 $Y=4350
XXFC9F1AD06 7 A<3> 5 WL<5> GND! VDD! 38 39 25 VDD! nor_5 $T=3238 3420 0 0 $X=2824 $Y=3202
XXFC9F1AD07 7 6 A<2> WL<6> GND! VDD! 40 41 26 VDD! nor_5 $T=3238 2272 0 0 $X=2824 $Y=2054
XXFC9F1AD08 7 6 5 WL<7> GND! VDD! 42 43 27 VDD! nor_5 $T=3238 1124 0 0 $X=2824 $Y=906
XXFC9F1AD09 A<2> 5 GND! VDD! VDD! VDD! inv_2 $T=2192 342 0 0 $X=1970 $Y=134
XXFC9F1AD010 A<3> 6 GND! VDD! VDD! VDD! inv_2 $T=1310 342 0 0 $X=1088 $Y=134
XXFC9F1AD011 A<4> 7 GND! VDD! VDD! VDD! inv_2 $T=460 342 0 0 $X=238 $Y=134
.ends rowdecoder
