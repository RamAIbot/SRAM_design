* PEX netlist file	Mon May  2 19:21:35 2022	tspc_flip_flop
* icv_netlist Version RHEL64 S-2021.06-SP2.6831572 2021/08/30
*.UNIT=4000

* Hierarchy Level 0

* Top of hierarchy  cell=tspc_flip_flop
.subckt tspc_flip_flop D 3 CLK 5 6 7 QBAR GND! VDD! 11 12
+	13
*.floating_nets _GENERATED_14 _GENERATED_15 _GENERATED_16 _GENERATED_17 _GENERATED_18 _GENERATED_19 _GENERATED_20 _GENERATED_21 _GENERATED_22 _GENERATED_23 _GENERATED_24
*+	_GENERATED_25 _GENERATED_26 _GENERATED_27
MM1 QBAR 7 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3458 $Y=1268  $PIN_XY=3488,1092,3458,1268,3428,1092 $DEVICE_ID=1001
MM2 7 6 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3122 $Y=1267  $PIN_XY=3152,1092,3122,1267,3092,1092 $DEVICE_ID=1001
MM3 6 CLK 13 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=2786 $Y=921  $PIN_XY=2816,922,2786,921,2756,922 $DEVICE_ID=1001
MM4 13 5 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=2618 $Y=914  $PIN_XY=2648,922,2618,914,2588,922 $DEVICE_ID=1001
MM5 5 3 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=2282 $Y=989  $PIN_XY=(2312,1092,2312,922),2282,989,(2252,1092,2252,922) $DEVICE_ID=1001
MM6 12 CLK GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=2114 $Y=1006  $PIN_XY=(2144,1092,2144,922),2114,1006,(2084,1092,2084,922) $DEVICE_ID=1001
MM7 3 D GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1778 $Y=920  $PIN_XY=1808,922,1778,920,1748,922 $DEVICE_ID=1001
MM8 QBAR 7 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3458 $Y=1268  $PIN_XY=(3488,1432,3488,1262),3458,1268,(3428,1432,3428,1262) $DEVICE_ID=1003
MM9 7 6 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3122 $Y=1267  $PIN_XY=(3152,1432,3152,1262),3122,1267,(3092,1432,3092,1262) $DEVICE_ID=1003
MM10 6 5 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2618 $Y=1455  $PIN_XY=2648,1432,2618,1455,2588,1432 $DEVICE_ID=1003
MM11 5 CLK VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2282 $Y=1452  $PIN_XY=2312,1432,2282,1452,2252,1432 $DEVICE_ID=1003
MM12 3 CLK 11 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=1946 $Y=1434  $PIN_XY=1976,1432,1946,1434,1916,1432 $DEVICE_ID=1003
MM13 11 D VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=1778 $Y=1434  $PIN_XY=1808,1432,1778,1434,1748,1432 $DEVICE_ID=1003
.ends tspc_flip_flop
