* PEX netlist file	Tue May  3 21:16:08 2022	bitcell
* icv_netlist Version RHEL64 S-2021.06-SP2.6831572 2021/08/30
*.UNIT=4000

* Hierarchy Level 0

* Top of hierarchy  cell=bitcell
.subckt bitcell 2 3 WL VDD! GND! BLB BL
*.floating_nets 5 6 11 12
MM1 BL WL 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=672 $Y=-164  $PIN_XY=702,-174,672,-164,642,-174 $DEVICE_ID=1001
MM2 GND! 2 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=336 $Y=-4  $PIN_XY=(366,0,366,-174),336,-4,(306,0,306,-174) $DEVICE_ID=1001
MM3 2 3 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=0 $Y=-4  $PIN_XY=(30,0,30,-174),0,-4,(-30,0,-30,-174) $DEVICE_ID=1001
MM4 2 WL BLB nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=-336 $Y=-164  $PIN_XY=-306,-174,-336,-164,-366,-174 $DEVICE_ID=1001
MM5 VDD! 2 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=336 $Y=-4  $PIN_XY=366,170,336,-4,306,170 $DEVICE_ID=1003
MM6 2 3 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=0 $Y=-4  $PIN_XY=30,170,0,-4,-30,170 $DEVICE_ID=1003
.ends bitcell
