* PEX netlist file	Wed May  4 03:42:47 2022	bit_cell_array
* icv_netlist Version RHEL64 S-2021.06-SP2.6831572 2021/08/30
*.UNIT=4000

* Hierarchy Level 3
.subckt bitcell 2 3 4 5 6 7 8 9 10 11 12
*.floating_nets _GENERATED_13
.ends bitcell
.subckt tspc_flip_flop 2 3 4 5 6 7 8 9 10 11 12
+	13 14 15
*.floating_nets _GENERATED_16 _GENERATED_17 _GENERATED_18 _GENERATED_19 _GENERATED_20 _GENERATED_21 _GENERATED_22 _GENERATED_23 _GENERATED_24 _GENERATED_25 _GENERATED_26
*+	_GENERATED_27
.ends tspc_flip_flop
.subckt inverter_write_driver 2 3 4 5 6 7 8 9 10
MM1 2 3 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=30 $Y=120  $PIN_XY=60,-76,30,120,0,-76 $DEVICE_ID=1001
MM2 2 3 8 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=30 $Y=120  $PIN_XY=60,316,30,120,0,316 $DEVICE_ID=1003
.ends inverter_write_driver
.subckt inv_2 2 3 4 5 6 7 8
.ends inv_2
.subckt nor_5 2 3 4 5 6 7 8 9 10 11
*.floating_nets _GENERATED_12 _GENERATED_13
.ends nor_5
.subckt and_2 2 3 4 5 6 7 8 9 10 11 12
*.floating_nets _GENERATED_13
MM1 5 3 6 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2450 $Y=1254  $PIN_XY=2480,1082,2450,1254,2420,1082 $DEVICE_ID=1001
.ends and_2

* Hierarchy Level 2
.subckt Write_Driver 3 4 6 7 18 19 20 21 22 23 24
*.floating_nets 14 15 16 17 _GENERATED_46 _GENERATED_47 _GENERATED_48 _GENERATED_49 _GENERATED_50 _GENERATED_51 _GENERATED_52
*+	_GENERATED_53
MM1 18 9 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1548 $Y=215  $PIN_XY=1578,252,1548,215,1518,252 $DEVICE_ID=1001
MM2 5 6 18 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1212 $Y=243  $PIN_XY=1242,252,1212,243,1182,252 $DEVICE_ID=1001
MM3 2 8 4 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=204 $Y=264  $PIN_XY=234,252,204,264,174,252 $DEVICE_ID=1001
MM4 5 8 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=-132 $Y=264  $PIN_XY=-102,252,-132,264,-162,252 $DEVICE_ID=1001
XX880FE34C36 9 6 10 _GENERATED_25 11 18 19 20 21 inverter_write_driver $T=846 328 0 0 $X=582 $Y=24
XX880FE34C37 8 7 12 13 10 18 19 20 21 inverter_write_driver $T=510 328 0 0 $X=246 $Y=24
.ends Write_Driver
.subckt bit_conditioning 3 4 5 6 7 8 9 10
*.floating_nets _GENERATED_19 _GENERATED_20 _GENERATED_21 _GENERATED_22
MM1 2 5 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3000 $Y=1838  $PIN_XY=3030,1668,3000,1838,2970,1668 $DEVICE_ID=1001
MM2 2 5 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3000 $Y=1838  $PIN_XY=(3030,2008,3030,1838),3000,1838,(2970,2008,2970,1838) $DEVICE_ID=1003
MM3 4 2 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2664 $Y=1838  $PIN_XY=2694,1838,2664,1838,2634,1838 $DEVICE_ID=1003
MM4 3 2 6 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2328 $Y=1838  $PIN_XY=2358,1838,2328,1838,2298,1838 $DEVICE_ID=1003
XX880FE34C38 5 2 7 6 8 9 10 inv_2 $T=3000 1668 0 0 $X=2778 $Y=1460
.ends bit_conditioning
.subckt rowdecoder 2 4 5 7 8 10 11 12 13 14 15
+	16 17
*.floating_nets 18 19 _GENERATED_159 _GENERATED_160 _GENERATED_161 _GENERATED_162 _GENERATED_163 _GENERATED_164 _GENERATED_165 _GENERATED_166 _GENERATED_167
*+	_GENERATED_168 _GENERATED_169 _GENERATED_170
MM1 10 2 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3722 $Y=9152  $PIN_XY=3752,9152,3722,9152,3692,9152 $DEVICE_ID=1001
MM2 11 2 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3722 $Y=8004  $PIN_XY=3752,8004,3722,8004,3692,8004 $DEVICE_ID=1001
MM3 12 3 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3722 $Y=6854  $PIN_XY=3752,6854,3722,6854,3692,6854 $DEVICE_ID=1001
MM4 13 3 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3722 $Y=5706  $PIN_XY=3752,5706,3722,5706,3692,5706 $DEVICE_ID=1001
MM5 14 2 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3722 $Y=4558  $PIN_XY=3752,4558,3722,4558,3692,4558 $DEVICE_ID=1001
MM6 15 2 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3722 $Y=3410  $PIN_XY=3752,3410,3722,3410,3692,3410 $DEVICE_ID=1001
MM7 16 3 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3722 $Y=2262  $PIN_XY=3752,2262,3722,2262,3692,2262 $DEVICE_ID=1001
MM8 17 3 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3722 $Y=1114  $PIN_XY=3752,1114,3722,1114,3692,1114 $DEVICE_ID=1001
MM9 10 8 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3386 $Y=9350  $PIN_XY=3416,9152,3386,9350,3356,9152 $DEVICE_ID=1001
MM10 11 9 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3386 $Y=8202  $PIN_XY=3416,8004,3386,8202,3356,8004 $DEVICE_ID=1001
MM11 12 8 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3386 $Y=7052  $PIN_XY=3416,6854,3386,7052,3356,6854 $DEVICE_ID=1001
MM12 13 9 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3386 $Y=5904  $PIN_XY=3416,5706,3386,5904,3356,5706 $DEVICE_ID=1001
MM13 14 8 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3386 $Y=4756  $PIN_XY=3416,4558,3386,4756,3356,4558 $DEVICE_ID=1001
MM14 15 9 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3386 $Y=3608  $PIN_XY=3416,3410,3386,3608,3356,3410 $DEVICE_ID=1001
MM15 16 8 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3386 $Y=2460  $PIN_XY=3416,2262,3386,2460,3356,2262 $DEVICE_ID=1001
MM16 17 9 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3386 $Y=1312  $PIN_XY=3416,1114,3386,1312,3356,1114 $DEVICE_ID=1001
MM17 10 5 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3050 $Y=9350  $PIN_XY=3080,9152,3050,9350,3020,9152 $DEVICE_ID=1001
MM18 11 5 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3050 $Y=8202  $PIN_XY=3080,8004,3050,8202,3020,8004 $DEVICE_ID=1001
MM19 12 5 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3050 $Y=7052  $PIN_XY=3080,6854,3050,7052,3020,6854 $DEVICE_ID=1001
MM20 13 5 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3050 $Y=5904  $PIN_XY=3080,5706,3050,5904,3020,5706 $DEVICE_ID=1001
MM21 14 6 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3050 $Y=4756  $PIN_XY=3080,4558,3050,4756,3020,4558 $DEVICE_ID=1001
MM22 15 6 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3050 $Y=3608  $PIN_XY=3080,3410,3050,3608,3020,3410 $DEVICE_ID=1001
MM23 16 6 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3050 $Y=2460  $PIN_XY=3080,2262,3050,2460,3020,2262 $DEVICE_ID=1001
MM24 17 6 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3050 $Y=1312  $PIN_XY=3080,1114,3050,1312,3020,1114 $DEVICE_ID=1001
MM25 9 8 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2192 $Y=512  $PIN_XY=2222,342,2192,512,2162,342 $DEVICE_ID=1001
MM26 3 2 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1310 $Y=512  $PIN_XY=1340,342,1310,512,1280,342 $DEVICE_ID=1001
MM27 6 5 7 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=460 $Y=512  $PIN_XY=490,342,460,512,430,342 $DEVICE_ID=1001
MM28 10 8 21 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3386 $Y=9350  $PIN_XY=(3416,9548,3416,9378),3386,9350,(3356,9548,3356,9378) $DEVICE_ID=1003
MM29 11 9 23 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3386 $Y=8202  $PIN_XY=(3416,8400,3416,8230),3386,8202,(3356,8400,3356,8230) $DEVICE_ID=1003
MM30 12 8 25 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3386 $Y=7052  $PIN_XY=(3416,7250,3416,7080),3386,7052,(3356,7250,3356,7080) $DEVICE_ID=1003
MM31 13 9 27 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3386 $Y=5904  $PIN_XY=(3416,6102,3416,5932),3386,5904,(3356,6102,3356,5932) $DEVICE_ID=1003
MM32 14 8 29 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3386 $Y=4756  $PIN_XY=(3416,4954,3416,4784),3386,4756,(3356,4954,3356,4784) $DEVICE_ID=1003
MM33 15 9 31 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3386 $Y=3608  $PIN_XY=(3416,3806,3416,3636),3386,3608,(3356,3806,3356,3636) $DEVICE_ID=1003
MM34 16 8 33 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3386 $Y=2460  $PIN_XY=(3416,2658,3416,2488),3386,2460,(3356,2658,3356,2488) $DEVICE_ID=1003
MM35 17 9 35 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3386 $Y=1312  $PIN_XY=(3416,1510,3416,1340),3386,1312,(3356,1510,3356,1340) $DEVICE_ID=1003
MM36 21 2 20 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=3218 $Y=9450  $PIN_XY=(3248,9548,3248,9378),3218,9450,(3188,9548,3188,9378) $DEVICE_ID=1003
MM37 23 2 22 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=3218 $Y=8302  $PIN_XY=(3248,8400,3248,8230),3218,8302,(3188,8400,3188,8230) $DEVICE_ID=1003
MM38 25 3 24 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=3218 $Y=7152  $PIN_XY=(3248,7250,3248,7080),3218,7152,(3188,7250,3188,7080) $DEVICE_ID=1003
MM39 27 3 26 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=3218 $Y=6004  $PIN_XY=(3248,6102,3248,5932),3218,6004,(3188,6102,3188,5932) $DEVICE_ID=1003
MM40 29 2 28 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=3218 $Y=4856  $PIN_XY=(3248,4954,3248,4784),3218,4856,(3188,4954,3188,4784) $DEVICE_ID=1003
MM41 31 2 30 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=3218 $Y=3708  $PIN_XY=(3248,3806,3248,3636),3218,3708,(3188,3806,3188,3636) $DEVICE_ID=1003
MM42 33 3 32 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=3218 $Y=2560  $PIN_XY=(3248,2658,3248,2488),3218,2560,(3188,2658,3188,2488) $DEVICE_ID=1003
MM43 35 3 34 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=1.134e-15 PDEO=2.34e-07
+	 PSEO=2.34e-07 $X=3218 $Y=1412  $PIN_XY=(3248,1510,3248,1340),3218,1412,(3188,1510,3188,1340) $DEVICE_ID=1003
MM44 20 5 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3050 $Y=9350  $PIN_XY=(3080,9548,3080,9378),3050,9350,(3020,9548,3020,9378) $DEVICE_ID=1003
MM45 22 5 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3050 $Y=8202  $PIN_XY=(3080,8400,3080,8230),3050,8202,(3020,8400,3020,8230) $DEVICE_ID=1003
MM46 24 5 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3050 $Y=7052  $PIN_XY=(3080,7250,3080,7080),3050,7052,(3020,7250,3020,7080) $DEVICE_ID=1003
MM47 26 5 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3050 $Y=5904  $PIN_XY=(3080,6102,3080,5932),3050,5904,(3020,6102,3020,5932) $DEVICE_ID=1003
MM48 28 6 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3050 $Y=4756  $PIN_XY=(3080,4954,3080,4784),3050,4756,(3020,4954,3020,4784) $DEVICE_ID=1003
MM49 30 6 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3050 $Y=3608  $PIN_XY=(3080,3806,3080,3636),3050,3608,(3020,3806,3020,3636) $DEVICE_ID=1003
MM50 32 6 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3050 $Y=2460  $PIN_XY=(3080,2658,3080,2488),3050,2460,(3020,2658,3020,2488) $DEVICE_ID=1003
MM51 34 6 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3050 $Y=1312  $PIN_XY=(3080,1510,3080,1340),3050,1312,(3020,1510,3020,1340) $DEVICE_ID=1003
MM52 9 8 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2192 $Y=512  $PIN_XY=(2222,682,2222,512),2192,512,(2162,682,2162,512) $DEVICE_ID=1003
MM53 3 2 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1310 $Y=512  $PIN_XY=(1340,682,1340,512),1310,512,(1280,682,1280,512) $DEVICE_ID=1003
MM54 6 5 4 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=460 $Y=512  $PIN_XY=(490,682,490,512),460,512,(430,682,430,512) $DEVICE_ID=1003
XX880FE34C39 2 5 8 10 7 4 20 21 4 36 nor_5 $T=3238 9162 0 0 $X=2824 $Y=8944
XX880FE34C40 2 5 9 11 7 4 22 23 4 37 nor_5 $T=3238 8014 0 0 $X=2824 $Y=7795
XX880FE34C41 3 5 8 12 7 4 24 25 4 38 nor_5 $T=3238 6864 0 0 $X=2824 $Y=6646
XX880FE34C42 3 5 9 13 7 4 26 27 4 39 nor_5 $T=3238 5716 0 0 $X=2824 $Y=5498
XX880FE34C43 2 6 8 14 7 4 28 29 4 40 nor_5 $T=3238 4568 0 0 $X=2824 $Y=4350
XX880FE34C44 2 6 9 15 7 4 30 31 4 41 nor_5 $T=3238 3420 0 0 $X=2824 $Y=3202
XX880FE34C45 3 6 8 16 7 4 32 33 4 42 nor_5 $T=3238 2272 0 0 $X=2824 $Y=2054
XX880FE34C46 3 6 9 17 7 4 34 35 4 43 nor_5 $T=3238 1124 0 0 $X=2824 $Y=906
XX880FE34C47 8 9 7 4 _GENERATED_44 4 4 inv_2 $T=2192 342 0 0 $X=1970 $Y=134
XX880FE34C48 2 3 7 4 _GENERATED_45 4 4 inv_2 $T=1310 342 0 0 $X=1088 $Y=134
XX880FE34C49 5 6 7 4 _GENERATED_46 4 4 inv_2 $T=460 342 0 0 $X=238 $Y=134
.ends rowdecoder
.subckt demu_2_4 4 5 6 7 8 9 10 15 17
*.floating_nets _GENERATED_89 _GENERATED_90 _GENERATED_91
MM1 13 4 23 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=3476 $Y=382  $PIN_XY=(3506,492,3506,322),3476,382,(3446,492,3446,322) $DEVICE_ID=1001
MM2 23 5 6 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=3308 $Y=577  $PIN_XY=(3338,492,3338,322),3308,577,(3278,492,3278,322) $DEVICE_ID=1001
MM3 12 3 21 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=2468 $Y=382  $PIN_XY=(2498,492,2498,322),2468,382,(2438,492,2438,322) $DEVICE_ID=1001
MM4 21 5 6 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=2300 $Y=577  $PIN_XY=(2330,492,2330,322),2300,577,(2270,492,2270,322) $DEVICE_ID=1001
MM5 11 4 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=1460 $Y=382  $PIN_XY=(1490,492,1490,322),1460,382,(1430,492,1430,322) $DEVICE_ID=1001
MM6 19 2 6 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=1292 $Y=577  $PIN_XY=(1322,492,1322,322),1292,577,(1262,492,1262,322) $DEVICE_ID=1001
MM7 6 5 2 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=620 $Y=1294  $PIN_XY=650,1462,620,1294,590,1462 $DEVICE_ID=1001
MM8 14 3 24 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=452 $Y=382  $PIN_XY=(482,492,482,322),452,382,(422,492,422,322) $DEVICE_ID=1001
MM9 6 4 3 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=284 $Y=1294  $PIN_XY=314,1462,284,1294,254,1462 $DEVICE_ID=1001
MM10 24 2 6 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=284 $Y=575  $PIN_XY=(314,492,314,322),284,575,(254,492,254,322) $DEVICE_ID=1001
MM11 9 13 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3980 $Y=664  $PIN_XY=(4010,832,4010,662),3980,664,(3950,832,3950,662) $DEVICE_ID=1003
MM12 13 4 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3644 $Y=765  $PIN_XY=(3674,832,3674,662),3644,765,(3614,832,3614,662) $DEVICE_ID=1003
MM13 13 5 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3308 $Y=577  $PIN_XY=(3338,832,3338,662),3308,577,(3278,832,3278,662) $DEVICE_ID=1003
MM14 8 12 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2972 $Y=664  $PIN_XY=(3002,832,3002,662),2972,664,(2942,832,2942,662) $DEVICE_ID=1003
MM15 12 3 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2636 $Y=765  $PIN_XY=(2666,832,2666,662),2636,765,(2606,832,2606,662) $DEVICE_ID=1003
MM16 12 5 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2300 $Y=577  $PIN_XY=(2330,832,2330,662),2300,577,(2270,832,2270,662) $DEVICE_ID=1003
MM17 7 11 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1964 $Y=664  $PIN_XY=(1994,832,1994,662),1964,664,(1934,832,1934,662) $DEVICE_ID=1003
MM18 11 4 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1628 $Y=765  $PIN_XY=(1658,832,1658,662),1628,765,(1598,832,1598,662) $DEVICE_ID=1003
MM19 11 2 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1292 $Y=577  $PIN_XY=(1322,832,1322,662),1292,577,(1262,832,1262,662) $DEVICE_ID=1003
MM20 10 14 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=956 $Y=664  $PIN_XY=(986,832,986,662),956,664,(926,832,926,662) $DEVICE_ID=1003
MM21 15 5 2 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=620 $Y=1294  $PIN_XY=(650,1292,650,1122),620,1294,(590,1292,590,1122) $DEVICE_ID=1003
MM22 14 3 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=620 $Y=763  $PIN_XY=(650,832,650,662),620,763,(590,832,590,662) $DEVICE_ID=1003
MM23 15 4 3 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=284 $Y=1294  $PIN_XY=(314,1292,314,1122),284,1294,(254,1292,254,1122) $DEVICE_ID=1003
MM24 14 2 15 pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=284 $Y=575  $PIN_XY=(314,832,314,662),284,575,(254,832,254,662) $DEVICE_ID=1003
XX880FE34C50 4 11 2 7 6 15 19 16 17 17 18 and_2 $T=-486 -590 0 0 $X=1070 $Y=113
XX880FE34C51 3 12 5 8 6 15 21 16 17 17 20 and_2 $T=522 -590 0 0 $X=2078 $Y=113
XX880FE34C52 4 13 5 9 6 15 23 16 17 17 22 and_2 $T=1530 -590 0 0 $X=3086 $Y=113
XX880FE34C53 3 14 2 10 6 15 24 16 17 17 6 and_2 $T=-1494 -590 0 0 $X=62 $Y=113
XX880FE34C54 5 2 6 15 16 17 17 inv_2 $T=620 1462 0 180 $X=398 $Y=913
XX880FE34C55 4 3 6 15 16 17 17 inv_2 $T=284 1462 0 180 $X=62 $Y=913
.ends demu_2_4
.subckt VCELLR4 2 3 4 5 6 7 8 9 10 11 12
+	13 14 15 16 17 18 19 20 21 22 23
+	24 25 26 27 28 29 30 31 32 33 34
+	35 36 37 38 39 40 41 42 43 44 45
+	46 47 48 49 50 51 52 53 54 55 56
+	57 58 59 60 61 62 63 64 65 66 67
+	68 69 70 71 72 73 74 75
*.floating_nets _GENERATED_172 _GENERATED_173 _GENERATED_174 _GENERATED_175 _GENERATED_176 _GENERATED_177 _GENERATED_178 _GENERATED_179 _GENERATED_180 _GENERATED_181 _GENERATED_182
*+	_GENERATED_183 _GENERATED_184 _GENERATED_185 _GENERATED_186 _GENERATED_187 _GENERATED_188 _GENERATED_189 _GENERATED_190 _GENERATED_191 _GENERATED_192
XX880FE34C58 11 10 2 26 27 44 43 58 59 74 75 bitcell $T=0 0 0 0 $X=-558 $Y=-410
XX880FE34C59 13 12 3 28 29 46 45 60 61 74 75 bitcell $T=1344 0 0 0 $X=786 $Y=-410
XX880FE34C60 15 14 4 30 31 48 47 62 63 74 75 bitcell $T=2688 0 0 0 $X=2130 $Y=-410
XX880FE34C61 17 16 5 32 33 50 49 64 65 74 75 bitcell $T=4032 0 0 0 $X=3474 $Y=-410
XX880FE34C62 19 18 6 34 35 42 51 66 67 74 75 bitcell $T=5376 0 0 0 $X=4818 $Y=-410
XX880FE34C63 21 20 7 36 37 53 52 68 69 74 75 bitcell $T=6720 0 0 0 $X=6162 $Y=-410
XX880FE34C64 23 22 8 38 39 55 54 70 71 74 75 bitcell $T=8064 0 0 0 $X=7506 $Y=-410
XX880FE34C65 25 24 9 40 41 57 56 72 73 74 75 bitcell $T=9408 0 0 0 $X=8850 $Y=-410
.ends VCELLR4

* Hierarchy Level 1
.subckt column_decoder_new 2 7 8 9 10 11 12 13 14 15 16
+	17 18 19 20 21 22 23 24 25 26 27
+	28 29 30 31 32 33 34 35 36 37 38
+	39 40 41 42 43 44 45 46 47 48 49
+	50
MM1 38 6 47 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10666 $Y=385  $PIN_XY=10696,380,10666,385,10636,380 $DEVICE_ID=1001
MM2 37 6 46 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10330 $Y=385  $PIN_XY=10360,380,10330,385,10300,380 $DEVICE_ID=1001
MM3 36 6 45 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9994 $Y=385  $PIN_XY=10024,380,9994,385,9964,380 $DEVICE_ID=1001
MM4 35 6 44 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9658 $Y=385  $PIN_XY=9688,380,9658,385,9628,380 $DEVICE_ID=1001
MM5 34 6 43 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9322 $Y=385  $PIN_XY=9352,380,9322,385,9292,380 $DEVICE_ID=1001
MM6 33 6 42 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8986 $Y=385  $PIN_XY=9016,380,8986,385,8956,380 $DEVICE_ID=1001
MM7 32 6 41 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8650 $Y=385  $PIN_XY=8680,380,8650,385,8620,380 $DEVICE_ID=1001
MM8 31 6 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8314 $Y=385  $PIN_XY=8344,380,8314,385,8284,380 $DEVICE_ID=1001
MM9 30 5 47 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7978 $Y=385  $PIN_XY=8008,380,7978,385,7948,380 $DEVICE_ID=1001
MM10 29 5 46 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7642 $Y=385  $PIN_XY=7672,380,7642,385,7612,380 $DEVICE_ID=1001
MM11 28 5 45 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7306 $Y=385  $PIN_XY=7336,380,7306,385,7276,380 $DEVICE_ID=1001
MM12 27 5 44 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6970 $Y=385  $PIN_XY=7000,380,6970,385,6940,380 $DEVICE_ID=1001
MM13 26 5 43 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6634 $Y=385  $PIN_XY=6664,380,6634,385,6604,380 $DEVICE_ID=1001
MM14 25 5 42 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6298 $Y=385  $PIN_XY=6328,380,6298,385,6268,380 $DEVICE_ID=1001
MM15 24 5 41 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5962 $Y=385  $PIN_XY=5992,380,5962,385,5932,380 $DEVICE_ID=1001
MM16 23 5 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5626 $Y=385  $PIN_XY=5656,380,5626,385,5596,380 $DEVICE_ID=1001
MM17 22 4 47 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5290 $Y=385  $PIN_XY=5320,380,5290,385,5260,380 $DEVICE_ID=1001
MM18 21 4 46 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4954 $Y=385  $PIN_XY=4984,380,4954,385,4924,380 $DEVICE_ID=1001
MM19 20 4 45 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4618 $Y=385  $PIN_XY=4648,380,4618,385,4588,380 $DEVICE_ID=1001
MM20 19 4 44 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4282 $Y=385  $PIN_XY=4312,380,4282,385,4252,380 $DEVICE_ID=1001
MM21 18 4 43 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3946 $Y=385  $PIN_XY=3976,380,3946,385,3916,380 $DEVICE_ID=1001
MM22 17 4 42 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3610 $Y=385  $PIN_XY=3640,380,3610,385,3580,380 $DEVICE_ID=1001
MM23 16 4 41 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3274 $Y=385  $PIN_XY=3304,380,3274,385,3244,380 $DEVICE_ID=1001
MM24 15 4 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2938 $Y=385  $PIN_XY=2968,380,2938,385,2908,380 $DEVICE_ID=1001
MM25 14 3 47 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2602 $Y=385  $PIN_XY=2632,380,2602,385,2572,380 $DEVICE_ID=1001
MM26 13 3 46 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2266 $Y=385  $PIN_XY=2296,380,2266,385,2236,380 $DEVICE_ID=1001
MM27 12 3 45 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1930 $Y=385  $PIN_XY=1960,380,1930,385,1900,380 $DEVICE_ID=1001
MM28 11 3 44 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1594 $Y=385  $PIN_XY=1624,380,1594,385,1564,380 $DEVICE_ID=1001
MM29 10 3 43 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1258 $Y=385  $PIN_XY=1288,380,1258,385,1228,380 $DEVICE_ID=1001
MM30 9 3 42 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=922 $Y=385  $PIN_XY=952,380,922,385,892,380 $DEVICE_ID=1001
MM31 8 3 41 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=586 $Y=385  $PIN_XY=616,380,586,385,556,380 $DEVICE_ID=1001
MM32 40 3 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=250 $Y=385  $PIN_XY=280,380,250,385,220,380 $DEVICE_ID=1001
XX880FE34C35 2 7 49 4 5 6 3 48 50 demu_2_4 $T=-6216 -556 0 0 $X=-6342 $Y=-442
.ends column_decoder_new
.subckt VCELLR2 2 3 4 5 6 7 8 9 10 11 12
+	13 14
XX880FE34C56 2 3 4 8 9 12 13 14 bit_conditioning $T=0 0 0 0 $X=2106 $Y=1348
XX880FE34C57 5 6 7 10 11 12 13 14 bit_conditioning $T=1008 0 0 0 $X=3114 $Y=1348
.ends VCELLR2

* Hierarchy Level 0

* Top of hierarchy  cell=bit_cell_array
.subckt bit_cell_array 2 3 4 5 6 7 8 9 VDD! GND! 12
+	13 CLK 15 16 17 18 19 20 21 22 23
+	24 25 26 27 28 29 30 31 32 33 34
+	35 36 37 38 39 40 41 42 43 44 WENB
+	D<0> D<1> D<3> D<2> A<4> A<3> A<2> 53 54 55 56
+	57 58 59 60 A<0> A<1> Q<3> Q<1> Q<0> Q<2>
*.floating_nets 595 596 597 598 599 600 601 602 603 604 605
*+	606 607 608 609 610 611 612 613 614 615 616
*+	617 618 619 620 621 622 623 624 625 626 627
*+	628 629 630 631 632 633 634 635 636 637 638
*+	639 640 641 642 643 644 645 646 647 648 649
*+	650 651 652 653 654 655 656 657 658 659 660
*+	661 662 663 664 665 666 667 668 669 670 671
*+	672 673 674 675 676 677 678 679 680 681 682
*+	683 684 685 686 687 688 689 690 691 692 693
*+	694 695 696 697 698 699 700 701 702 703 704
*+	705 706 707 708 709 710 711 712 713 714 715
*+	716 717 718 719 720 721 722 723 724 725 726
*+	727 728 729 730 731 732 733 734 735 736 737
*+	738 739 740 741 742 743 744 745 746 747 748
*+	749 750 751 752 753 754 755 756 757 758 759
*+	760 761 762 763 764 765 766 767 768 769 770
*+	771 772 773 774 775 776 777 778 779 780 781
*+	782 783 784 785 786 787 788 789 790 791 792
*+	793 794 795 796 797 798 799 800 801 802 803
*+	804 805 806 807 808 809 810 811 812 813 814
*+	815 816 817 818 819 820 821 822 823 824 825
*+	826 827 828 829 830 831 832 833 834 835 836
*+	837 838 839 840 841 842 843 844 845 846 847
*+	848 849 850 851 852 853 854 855 856 857 858
*+	859 860 861 862 863 864 865 866 867 868 869
*+	870 871 872 873 874 875 876 877 878 879 880
*+	881 882 883 884 885 886 887 888 889 890 891
*+	892 893 894 895 896 897 898 899 900 901 902
*+	903 904 905 906 907 908 909 910 911 912 913
*+	914 915 916 917 918 919 920 921 922 923 924
*+	925 926 927 928 929 930 931 932 933 934 935
*+	936 937 938 939 940 941 942 943 944 945 946
*+	947 948 949 950 951 952 953 954 955 956 957
*+	958 959 960 961 962 963 964 965 966 967 968
*+	969 970 971 972 973 974 975 976 977 978 979
*+	980 981 982 983 984 985 986 987 988 989 990
*+	991 992 993 994 995 996 997 998 999 1000 1001
*+	1002 1003 1004 1005 1006 1007 1008 1009 1010 1011 1012
*+	1013 1014 1015 1016 1017 1018 1019 1020 1021 1022 1023
*+	1024 1025 1026 1027 1028 1029 1030 1031 1032 1033 1034
*+	1035 1036 1037 1038 1039 1040 1041 1042 1043 1044 1045
*+	1046 1047 1048 1049 1050 1051 1052 1053 1054 1055 1056
*+	1057 1058 1059 1060 1061 1062 1063 1064 1065 1066 1067
*+	1068 1069 1070 1071 1072 1073 1074 1075 1076 1077 1078
*+	1079 1080 1081 1082 1083 1084 1085 1086 1087 1088 1089
*+	1090 1091 1092 1093 1094 1095 1096 1097 1098 1099 1100
*+	1101 1102 1103 1104 1105 1106 1107 1108 1109 1110 1111
*+	1112 1113 1114 1115 1116 1117 1118 1119 1120 1121 1122
*+	1123 1124 1125 1126 1127 1128 1129 1130 1131 1132 1133
*+	1134 1135 1136 1137 1138 1139 1140 1141 1142 1143 1144
*+	1145 1146 1147 1148 1149 1150 1151 1152 1153 1154 1155
*+	1156 1157 1158 1159 1160 1161 1162 1163 1164 1165 1166
*+	1167 1168 1169 1170 1171 1172 1173 1174 1175 1176 1177
*+	1178 1179 1180 1181 1182 1183 1184 1185 1186 1187 1188
*+	1189 1190 1191 1192 1193 1194 1195 1196 1197 1198 1199
*+	1200 1201 1202 1203 1204 1205 1206 1207 1208 1209 1210
*+	1211 1212 1213 1214 1215 1216 1217 1218 1219 1220 1221
*+	1222 1223 1224 1225 1226 1227 1228 1229 1230 1231 1232
*+	1233 1234 1235 1236 1237 1238 1239 1240 1241 1242 1243
*+	1244 1245 1246 1247 1248 1249 1250 1251 1252 1253 1254
*+	1255 1256 1257 1258 1259 1260 1261 1262 1263 1264 1265
*+	1266 1267 1268 1269 1270 1271 1272 1273 1274 1275 1276
*+	1277 1278 1279 1280 1281 1282 1283 1284 1285 1286 1287
*+	1288 1289 1290 1291 1292 1293 1294 1295 1296 1297 1298
*+	1299 1300 1301 1302 1303 1304 1305 1306 1307 1308 1309
*+	1310 1311 1312 1313 1314 1315 1316 1317 1318 1319 1320
*+	1321 1322 1323 1324 1325 1326 1327 1328 1329 1330 1331
*+	1332 1333 1334 1335 1336 1337 1338 1339 1340 1341 1342
*+	1343 1344 1345 1346 1347 1348 1349 1350 1351 1352 1353
*+	1354 1355 1356 1357 1358 1359 1360 1361 1362 1363 1364
*+	1365 1366 1367 1368 1369 1370 1371 1372 1373 1374 1375
*+	1376 1377 1378 1379 1380 1381 1382 1383 1384 1385 1386
*+	1387 1388 1389 1390 1391 1392 1393 1394 1395 1396 1397
*+	1398 1399 1400 1401 1402 1403 1404 1405 1406 1407 1408
*+	1409 1410 1411 1412 1413 1414 1415 1416 1417 1418 1419
*+	1420 1421 1422 1423 1424 1425 1426 1427 1428 1429 1430
*+	1431 1432 1433 1434 1435 1436 1437 1438 1439 1440 1441
*+	1442 1443 1444 1445 1446 1447 1448 1449 1450 1451 1452
*+	1453 1454 1455 1456 1457 1458 1459 1460 1461 1462 1463
*+	1464 1465 1466 1467 1468 1469 1470 1471 1472 1473 1474
*+	1475 1476 1477 1478 1479 1480 1481 1482 1483 1484 1485
*+	1486 1487 1488 1489 1490 1491 1492 1493 1494 1495 1496
*+	1497 1498 1499 1500 1501 1502 1503 1504 1505 1506 1507
*+	1508 1509 1510 1511 1512 1513 1514 1515 1516 1517 1518
*+	1519 1520 _GENERATED_5219 _GENERATED_5220 _GENERATED_5221 _GENERATED_5222 _GENERATED_5223 _GENERATED_5224 _GENERATED_5225 _GENERATED_5226 _GENERATED_5227
*+	_GENERATED_5228 _GENERATED_5229 _GENERATED_5230 _GENERATED_5231 _GENERATED_5232 _GENERATED_5233 _GENERATED_5234 _GENERATED_5235 _GENERATED_5236 _GENERATED_5237 _GENERATED_5238
*+	_GENERATED_5239 _GENERATED_5240 _GENERATED_5241 _GENERATED_5242 _GENERATED_5243 _GENERATED_5244 _GENERATED_5245 _GENERATED_5246 _GENERATED_5247 _GENERATED_5248 _GENERATED_5249
MM1 44 60 321 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20676 $Y=75  $PIN_XY=20706,158,20676,75,20646,158 $DEVICE_ID=1001
MM2 44 59 289 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20676 $Y=-1072  $PIN_XY=20706,-990,20676,-1072,20646,-990 $DEVICE_ID=1001
MM3 44 58 257 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20676 $Y=-2219  $PIN_XY=20706,-2136,20676,-2219,20646,-2136 $DEVICE_ID=1001
MM4 GND! 322 321 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=20340 $Y=304  $PIN_XY=(20370,332,20370,158),20340,304,(20310,332,20310,158) $DEVICE_ID=1001
MM5 GND! 290 289 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=20340 $Y=-720  $PIN_XY=(20370,-816,20370,-990),20340,-720,(20310,-816,20310,-990) $DEVICE_ID=1001
MM6 GND! 258 257 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=20340 $Y=-1867  $PIN_XY=(20370,-1962,20370,-2136),20340,-1867,(20310,-1962,20310,-2136) $DEVICE_ID=1001
MM7 322 321 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=20004 $Y=304  $PIN_XY=(20034,332,20034,158),20004,304,(19974,332,19974,158) $DEVICE_ID=1001
MM8 290 289 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=20004 $Y=-720  $PIN_XY=(20034,-816,20034,-990),20004,-720,(19974,-816,19974,-990) $DEVICE_ID=1001
MM9 258 257 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=20004 $Y=-1867  $PIN_XY=(20034,-1962,20034,-2136),20004,-1867,(19974,-1962,19974,-2136) $DEVICE_ID=1001
MM10 322 60 43 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=19668 $Y=75  $PIN_XY=19698,158,19668,75,19638,158 $DEVICE_ID=1001
MM11 290 59 43 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=19668 $Y=-1072  $PIN_XY=19698,-990,19668,-1072,19638,-990 $DEVICE_ID=1001
MM12 258 58 43 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=19668 $Y=-2219  $PIN_XY=19698,-2136,19668,-2219,19638,-2136 $DEVICE_ID=1001
MM13 42 60 319 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=19332 $Y=75  $PIN_XY=19362,158,19332,75,19302,158 $DEVICE_ID=1001
MM14 42 59 287 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=19332 $Y=-1072  $PIN_XY=19362,-990,19332,-1072,19302,-990 $DEVICE_ID=1001
MM15 42 58 255 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=19332 $Y=-2219  $PIN_XY=19362,-2136,19332,-2219,19302,-2136 $DEVICE_ID=1001
MM16 GND! 320 319 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=18996 $Y=304  $PIN_XY=(19026,332,19026,158),18996,304,(18966,332,18966,158) $DEVICE_ID=1001
MM17 GND! 288 287 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=18996 $Y=-720  $PIN_XY=(19026,-816,19026,-990),18996,-720,(18966,-816,18966,-990) $DEVICE_ID=1001
MM18 GND! 256 255 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=18996 $Y=-1867  $PIN_XY=(19026,-1962,19026,-2136),18996,-1867,(18966,-1962,18966,-2136) $DEVICE_ID=1001
MM19 320 319 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=18660 $Y=304  $PIN_XY=(18690,332,18690,158),18660,304,(18630,332,18630,158) $DEVICE_ID=1001
MM20 288 287 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=18660 $Y=-720  $PIN_XY=(18690,-816,18690,-990),18660,-720,(18630,-816,18630,-990) $DEVICE_ID=1001
MM21 256 255 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=18660 $Y=-1867  $PIN_XY=(18690,-1962,18690,-2136),18660,-1867,(18630,-1962,18630,-2136) $DEVICE_ID=1001
MM22 320 60 41 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18324 $Y=75  $PIN_XY=18354,158,18324,75,18294,158 $DEVICE_ID=1001
MM23 288 59 41 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18324 $Y=-1072  $PIN_XY=18354,-990,18324,-1072,18294,-990 $DEVICE_ID=1001
MM24 256 58 41 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18324 $Y=-2219  $PIN_XY=18354,-2136,18324,-2219,18294,-2136 $DEVICE_ID=1001
MM25 40 60 317 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17988 $Y=75  $PIN_XY=18018,158,17988,75,17958,158 $DEVICE_ID=1001
MM26 40 59 285 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17988 $Y=-1072  $PIN_XY=18018,-990,17988,-1072,17958,-990 $DEVICE_ID=1001
MM27 40 58 253 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17988 $Y=-2219  $PIN_XY=18018,-2136,17988,-2219,17958,-2136 $DEVICE_ID=1001
MM28 GND! 318 317 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17652 $Y=304  $PIN_XY=(17682,332,17682,158),17652,304,(17622,332,17622,158) $DEVICE_ID=1001
MM29 GND! 286 285 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17652 $Y=-720  $PIN_XY=(17682,-816,17682,-990),17652,-720,(17622,-816,17622,-990) $DEVICE_ID=1001
MM30 GND! 254 253 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17652 $Y=-1867  $PIN_XY=(17682,-1962,17682,-2136),17652,-1867,(17622,-1962,17622,-2136) $DEVICE_ID=1001
MM31 318 317 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17316 $Y=304  $PIN_XY=(17346,332,17346,158),17316,304,(17286,332,17286,158) $DEVICE_ID=1001
MM32 286 285 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17316 $Y=-720  $PIN_XY=(17346,-816,17346,-990),17316,-720,(17286,-816,17286,-990) $DEVICE_ID=1001
MM33 254 253 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17316 $Y=-1867  $PIN_XY=(17346,-1962,17346,-2136),17316,-1867,(17286,-1962,17286,-2136) $DEVICE_ID=1001
MM34 318 60 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16980 $Y=75  $PIN_XY=17010,158,16980,75,16950,158 $DEVICE_ID=1001
MM35 286 59 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16980 $Y=-1072  $PIN_XY=17010,-990,16980,-1072,16950,-990 $DEVICE_ID=1001
MM36 254 58 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16980 $Y=-2219  $PIN_XY=17010,-2136,16980,-2219,16950,-2136 $DEVICE_ID=1001
MM37 38 60 315 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16644 $Y=75  $PIN_XY=16674,158,16644,75,16614,158 $DEVICE_ID=1001
MM38 38 59 283 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16644 $Y=-1072  $PIN_XY=16674,-990,16644,-1072,16614,-990 $DEVICE_ID=1001
MM39 38 58 251 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16644 $Y=-2219  $PIN_XY=16674,-2136,16644,-2219,16614,-2136 $DEVICE_ID=1001
MM40 GND! 316 315 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=16308 $Y=304  $PIN_XY=(16338,332,16338,158),16308,304,(16278,332,16278,158) $DEVICE_ID=1001
MM41 GND! 284 283 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=16308 $Y=-720  $PIN_XY=(16338,-816,16338,-990),16308,-720,(16278,-816,16278,-990) $DEVICE_ID=1001
MM42 GND! 252 251 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=16308 $Y=-1867  $PIN_XY=(16338,-1962,16338,-2136),16308,-1867,(16278,-1962,16278,-2136) $DEVICE_ID=1001
MM43 316 315 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=15972 $Y=304  $PIN_XY=(16002,332,16002,158),15972,304,(15942,332,15942,158) $DEVICE_ID=1001
MM44 284 283 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=15972 $Y=-720  $PIN_XY=(16002,-816,16002,-990),15972,-720,(15942,-816,15942,-990) $DEVICE_ID=1001
MM45 252 251 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=15972 $Y=-1867  $PIN_XY=(16002,-1962,16002,-2136),15972,-1867,(15942,-1962,15942,-2136) $DEVICE_ID=1001
MM46 316 60 37 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15636 $Y=75  $PIN_XY=15666,158,15636,75,15606,158 $DEVICE_ID=1001
MM47 284 59 37 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15636 $Y=-1072  $PIN_XY=15666,-990,15636,-1072,15606,-990 $DEVICE_ID=1001
MM48 252 58 37 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15636 $Y=-2219  $PIN_XY=15666,-2136,15636,-2219,15606,-2136 $DEVICE_ID=1001
MM49 36 60 313 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15300 $Y=75  $PIN_XY=15330,158,15300,75,15270,158 $DEVICE_ID=1001
MM50 36 59 281 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15300 $Y=-1072  $PIN_XY=15330,-990,15300,-1072,15270,-990 $DEVICE_ID=1001
MM51 36 58 249 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15300 $Y=-2219  $PIN_XY=15330,-2136,15300,-2219,15270,-2136 $DEVICE_ID=1001
MM52 GND! 314 313 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14964 $Y=304  $PIN_XY=(14994,332,14994,158),14964,304,(14934,332,14934,158) $DEVICE_ID=1001
MM53 GND! 282 281 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14964 $Y=-720  $PIN_XY=(14994,-816,14994,-990),14964,-720,(14934,-816,14934,-990) $DEVICE_ID=1001
MM54 GND! 250 249 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14964 $Y=-1867  $PIN_XY=(14994,-1962,14994,-2136),14964,-1867,(14934,-1962,14934,-2136) $DEVICE_ID=1001
MM55 314 313 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14628 $Y=304  $PIN_XY=(14658,332,14658,158),14628,304,(14598,332,14598,158) $DEVICE_ID=1001
MM56 282 281 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14628 $Y=-720  $PIN_XY=(14658,-816,14658,-990),14628,-720,(14598,-816,14598,-990) $DEVICE_ID=1001
MM57 314 60 35 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14292 $Y=75  $PIN_XY=14322,158,14292,75,14262,158 $DEVICE_ID=1001
MM58 282 59 35 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14292 $Y=-1072  $PIN_XY=14322,-990,14292,-1072,14262,-990 $DEVICE_ID=1001
MM59 34 60 311 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13956 $Y=75  $PIN_XY=13986,158,13956,75,13926,158 $DEVICE_ID=1001
MM60 34 59 279 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13956 $Y=-1072  $PIN_XY=13986,-990,13956,-1072,13926,-990 $DEVICE_ID=1001
MM61 GND! 312 311 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13620 $Y=304  $PIN_XY=(13650,332,13650,158),13620,304,(13590,332,13590,158) $DEVICE_ID=1001
MM62 GND! 280 279 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13620 $Y=-720  $PIN_XY=(13650,-816,13650,-990),13620,-720,(13590,-816,13590,-990) $DEVICE_ID=1001
MM63 312 311 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13284 $Y=304  $PIN_XY=(13314,332,13314,158),13284,304,(13254,332,13254,158) $DEVICE_ID=1001
MM64 280 279 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13284 $Y=-720  $PIN_XY=(13314,-816,13314,-990),13284,-720,(13254,-816,13254,-990) $DEVICE_ID=1001
MM65 312 60 33 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12948 $Y=75  $PIN_XY=12978,158,12948,75,12918,158 $DEVICE_ID=1001
MM66 280 59 33 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12948 $Y=-1072  $PIN_XY=12978,-990,12948,-1072,12918,-990 $DEVICE_ID=1001
MM67 250 249 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14628 $Y=-1867  $PIN_XY=(14658,-1962,14658,-2136),14628,-1867,(14598,-1962,14598,-2136) $DEVICE_ID=1001
MM68 250 58 35 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14292 $Y=-2219  $PIN_XY=14322,-2136,14292,-2219,14262,-2136 $DEVICE_ID=1001
MM69 34 58 247 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13956 $Y=-2219  $PIN_XY=13986,-2136,13956,-2219,13926,-2136 $DEVICE_ID=1001
MM70 GND! 248 247 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13620 $Y=-1867  $PIN_XY=(13650,-1962,13650,-2136),13620,-1867,(13590,-1962,13590,-2136) $DEVICE_ID=1001
MM71 248 247 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13284 $Y=-1867  $PIN_XY=(13314,-1962,13314,-2136),13284,-1867,(13254,-1962,13254,-2136) $DEVICE_ID=1001
MM72 248 58 33 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12948 $Y=-2219  $PIN_XY=12978,-2136,12948,-2219,12918,-2136 $DEVICE_ID=1001
MM73 32 60 309 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12612 $Y=75  $PIN_XY=12642,158,12612,75,12582,158 $DEVICE_ID=1001
MM74 32 59 277 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12612 $Y=-1072  $PIN_XY=12642,-990,12612,-1072,12582,-990 $DEVICE_ID=1001
MM75 32 58 245 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12612 $Y=-2219  $PIN_XY=12642,-2136,12612,-2219,12582,-2136 $DEVICE_ID=1001
MM76 GND! 310 309 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=12276 $Y=304  $PIN_XY=(12306,332,12306,158),12276,304,(12246,332,12246,158) $DEVICE_ID=1001
MM77 GND! 278 277 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=12276 $Y=-720  $PIN_XY=(12306,-816,12306,-990),12276,-720,(12246,-816,12246,-990) $DEVICE_ID=1001
MM78 GND! 246 245 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=12276 $Y=-1867  $PIN_XY=(12306,-1962,12306,-2136),12276,-1867,(12246,-1962,12246,-2136) $DEVICE_ID=1001
MM79 310 309 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11940 $Y=304  $PIN_XY=(11970,332,11970,158),11940,304,(11910,332,11910,158) $DEVICE_ID=1001
MM80 278 277 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11940 $Y=-720  $PIN_XY=(11970,-816,11970,-990),11940,-720,(11910,-816,11910,-990) $DEVICE_ID=1001
MM81 246 245 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11940 $Y=-1867  $PIN_XY=(11970,-1962,11970,-2136),11940,-1867,(11910,-1962,11910,-2136) $DEVICE_ID=1001
MM82 310 60 31 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11604 $Y=75  $PIN_XY=11634,158,11604,75,11574,158 $DEVICE_ID=1001
MM83 278 59 31 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11604 $Y=-1072  $PIN_XY=11634,-990,11604,-1072,11574,-990 $DEVICE_ID=1001
MM84 246 58 31 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11604 $Y=-2219  $PIN_XY=11634,-2136,11604,-2219,11574,-2136 $DEVICE_ID=1001
MM85 30 60 307 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11268 $Y=75  $PIN_XY=11298,158,11268,75,11238,158 $DEVICE_ID=1001
MM86 30 59 275 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11268 $Y=-1072  $PIN_XY=11298,-990,11268,-1072,11238,-990 $DEVICE_ID=1001
MM87 30 58 243 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11268 $Y=-2219  $PIN_XY=11298,-2136,11268,-2219,11238,-2136 $DEVICE_ID=1001
MM88 GND! 308 307 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10932 $Y=304  $PIN_XY=(10962,332,10962,158),10932,304,(10902,332,10902,158) $DEVICE_ID=1001
MM89 GND! 276 275 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10932 $Y=-720  $PIN_XY=(10962,-816,10962,-990),10932,-720,(10902,-816,10902,-990) $DEVICE_ID=1001
MM90 GND! 244 243 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10932 $Y=-1867  $PIN_XY=(10962,-1962,10962,-2136),10932,-1867,(10902,-1962,10902,-2136) $DEVICE_ID=1001
MM91 308 307 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10596 $Y=304  $PIN_XY=(10626,332,10626,158),10596,304,(10566,332,10566,158) $DEVICE_ID=1001
MM92 308 60 29 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10260 $Y=75  $PIN_XY=10290,158,10260,75,10230,158 $DEVICE_ID=1001
MM93 28 60 305 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9924 $Y=75  $PIN_XY=9954,158,9924,75,9894,158 $DEVICE_ID=1001
MM94 GND! 306 305 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9588 $Y=304  $PIN_XY=(9618,332,9618,158),9588,304,(9558,332,9558,158) $DEVICE_ID=1001
MM95 306 305 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9252 $Y=304  $PIN_XY=(9282,332,9282,158),9252,304,(9222,332,9222,158) $DEVICE_ID=1001
MM96 306 60 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8916 $Y=75  $PIN_XY=8946,158,8916,75,8886,158 $DEVICE_ID=1001
MM97 276 275 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10596 $Y=-720  $PIN_XY=(10626,-816,10626,-990),10596,-720,(10566,-816,10566,-990) $DEVICE_ID=1001
MM98 244 243 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10596 $Y=-1867  $PIN_XY=(10626,-1962,10626,-2136),10596,-1867,(10566,-1962,10566,-2136) $DEVICE_ID=1001
MM99 276 59 29 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10260 $Y=-1072  $PIN_XY=10290,-990,10260,-1072,10230,-990 $DEVICE_ID=1001
MM100 244 58 29 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10260 $Y=-2219  $PIN_XY=10290,-2136,10260,-2219,10230,-2136 $DEVICE_ID=1001
MM101 28 59 273 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9924 $Y=-1072  $PIN_XY=9954,-990,9924,-1072,9894,-990 $DEVICE_ID=1001
MM102 28 58 241 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9924 $Y=-2219  $PIN_XY=9954,-2136,9924,-2219,9894,-2136 $DEVICE_ID=1001
MM103 GND! 274 273 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9588 $Y=-720  $PIN_XY=(9618,-816,9618,-990),9588,-720,(9558,-816,9558,-990) $DEVICE_ID=1001
MM104 GND! 242 241 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9588 $Y=-1867  $PIN_XY=(9618,-1962,9618,-2136),9588,-1867,(9558,-1962,9558,-2136) $DEVICE_ID=1001
MM105 274 273 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9252 $Y=-720  $PIN_XY=(9282,-816,9282,-990),9252,-720,(9222,-816,9222,-990) $DEVICE_ID=1001
MM106 242 241 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9252 $Y=-1867  $PIN_XY=(9282,-1962,9282,-2136),9252,-1867,(9222,-1962,9222,-2136) $DEVICE_ID=1001
MM107 274 59 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8916 $Y=-1072  $PIN_XY=8946,-990,8916,-1072,8886,-990 $DEVICE_ID=1001
MM108 242 58 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8916 $Y=-2219  $PIN_XY=8946,-2136,8916,-2219,8886,-2136 $DEVICE_ID=1001
MM109 26 60 303 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8580 $Y=75  $PIN_XY=8610,158,8580,75,8550,158 $DEVICE_ID=1001
MM110 26 59 271 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8580 $Y=-1072  $PIN_XY=8610,-990,8580,-1072,8550,-990 $DEVICE_ID=1001
MM111 GND! 304 303 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8244 $Y=304  $PIN_XY=(8274,332,8274,158),8244,304,(8214,332,8214,158) $DEVICE_ID=1001
MM112 GND! 272 271 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8244 $Y=-720  $PIN_XY=(8274,-816,8274,-990),8244,-720,(8214,-816,8214,-990) $DEVICE_ID=1001
MM113 304 303 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7908 $Y=304  $PIN_XY=(7938,332,7938,158),7908,304,(7878,332,7878,158) $DEVICE_ID=1001
MM114 272 271 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7908 $Y=-720  $PIN_XY=(7938,-816,7938,-990),7908,-720,(7878,-816,7878,-990) $DEVICE_ID=1001
MM115 304 60 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7572 $Y=75  $PIN_XY=7602,158,7572,75,7542,158 $DEVICE_ID=1001
MM116 272 59 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7572 $Y=-1072  $PIN_XY=7602,-990,7572,-1072,7542,-990 $DEVICE_ID=1001
MM117 24 60 301 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7236 $Y=75  $PIN_XY=7266,158,7236,75,7206,158 $DEVICE_ID=1001
MM118 24 59 269 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7236 $Y=-1072  $PIN_XY=7266,-990,7236,-1072,7206,-990 $DEVICE_ID=1001
MM119 GND! 302 301 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6900 $Y=304  $PIN_XY=(6930,332,6930,158),6900,304,(6870,332,6870,158) $DEVICE_ID=1001
MM120 GND! 270 269 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6900 $Y=-720  $PIN_XY=(6930,-816,6930,-990),6900,-720,(6870,-816,6870,-990) $DEVICE_ID=1001
MM121 26 58 239 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8580 $Y=-2219  $PIN_XY=8610,-2136,8580,-2219,8550,-2136 $DEVICE_ID=1001
MM122 GND! 240 239 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8244 $Y=-1867  $PIN_XY=(8274,-1962,8274,-2136),8244,-1867,(8214,-1962,8214,-2136) $DEVICE_ID=1001
MM123 240 239 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7908 $Y=-1867  $PIN_XY=(7938,-1962,7938,-2136),7908,-1867,(7878,-1962,7878,-2136) $DEVICE_ID=1001
MM124 240 58 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7572 $Y=-2219  $PIN_XY=7602,-2136,7572,-2219,7542,-2136 $DEVICE_ID=1001
MM125 24 58 237 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7236 $Y=-2219  $PIN_XY=7266,-2136,7236,-2219,7206,-2136 $DEVICE_ID=1001
MM126 GND! 238 237 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6900 $Y=-1867  $PIN_XY=(6930,-1962,6930,-2136),6900,-1867,(6870,-1962,6870,-2136) $DEVICE_ID=1001
MM127 302 301 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6564 $Y=304  $PIN_XY=(6594,332,6594,158),6564,304,(6534,332,6534,158) $DEVICE_ID=1001
MM128 270 269 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6564 $Y=-720  $PIN_XY=(6594,-816,6594,-990),6564,-720,(6534,-816,6534,-990) $DEVICE_ID=1001
MM129 238 237 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6564 $Y=-1867  $PIN_XY=(6594,-1962,6594,-2136),6564,-1867,(6534,-1962,6534,-2136) $DEVICE_ID=1001
MM130 302 60 23 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6228 $Y=75  $PIN_XY=6258,158,6228,75,6198,158 $DEVICE_ID=1001
MM131 270 59 23 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6228 $Y=-1072  $PIN_XY=6258,-990,6228,-1072,6198,-990 $DEVICE_ID=1001
MM132 238 58 23 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6228 $Y=-2219  $PIN_XY=6258,-2136,6228,-2219,6198,-2136 $DEVICE_ID=1001
MM133 22 60 299 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5892 $Y=75  $PIN_XY=5922,158,5892,75,5862,158 $DEVICE_ID=1001
MM134 22 59 267 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5892 $Y=-1072  $PIN_XY=5922,-990,5892,-1072,5862,-990 $DEVICE_ID=1001
MM135 22 58 235 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5892 $Y=-2219  $PIN_XY=5922,-2136,5892,-2219,5862,-2136 $DEVICE_ID=1001
MM136 GND! 300 299 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5556 $Y=304  $PIN_XY=(5586,332,5586,158),5556,304,(5526,332,5526,158) $DEVICE_ID=1001
MM137 GND! 268 267 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5556 $Y=-720  $PIN_XY=(5586,-816,5586,-990),5556,-720,(5526,-816,5526,-990) $DEVICE_ID=1001
MM138 GND! 236 235 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5556 $Y=-1867  $PIN_XY=(5586,-1962,5586,-2136),5556,-1867,(5526,-1962,5526,-2136) $DEVICE_ID=1001
MM139 300 299 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5220 $Y=304  $PIN_XY=(5250,332,5250,158),5220,304,(5190,332,5190,158) $DEVICE_ID=1001
MM140 268 267 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5220 $Y=-720  $PIN_XY=(5250,-816,5250,-990),5220,-720,(5190,-816,5190,-990) $DEVICE_ID=1001
MM141 236 235 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5220 $Y=-1867  $PIN_XY=(5250,-1962,5250,-2136),5220,-1867,(5190,-1962,5190,-2136) $DEVICE_ID=1001
MM142 300 60 21 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4884 $Y=75  $PIN_XY=4914,158,4884,75,4854,158 $DEVICE_ID=1001
MM143 268 59 21 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4884 $Y=-1072  $PIN_XY=4914,-990,4884,-1072,4854,-990 $DEVICE_ID=1001
MM144 236 58 21 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4884 $Y=-2219  $PIN_XY=4914,-2136,4884,-2219,4854,-2136 $DEVICE_ID=1001
MM145 20 60 297 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4548 $Y=75  $PIN_XY=4578,158,4548,75,4518,158 $DEVICE_ID=1001
MM146 20 59 265 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4548 $Y=-1072  $PIN_XY=4578,-990,4548,-1072,4518,-990 $DEVICE_ID=1001
MM147 20 58 233 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4548 $Y=-2219  $PIN_XY=4578,-2136,4548,-2219,4518,-2136 $DEVICE_ID=1001
MM148 GND! 298 297 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4212 $Y=304  $PIN_XY=(4242,332,4242,158),4212,304,(4182,332,4182,158) $DEVICE_ID=1001
MM149 GND! 266 265 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4212 $Y=-720  $PIN_XY=(4242,-816,4242,-990),4212,-720,(4182,-816,4182,-990) $DEVICE_ID=1001
MM150 GND! 234 233 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4212 $Y=-1867  $PIN_XY=(4242,-1962,4242,-2136),4212,-1867,(4182,-1962,4182,-2136) $DEVICE_ID=1001
MM151 298 297 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3876 $Y=304  $PIN_XY=(3906,332,3906,158),3876,304,(3846,332,3846,158) $DEVICE_ID=1001
MM152 266 265 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3876 $Y=-720  $PIN_XY=(3906,-816,3906,-990),3876,-720,(3846,-816,3846,-990) $DEVICE_ID=1001
MM153 234 233 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3876 $Y=-1867  $PIN_XY=(3906,-1962,3906,-2136),3876,-1867,(3846,-1962,3846,-2136) $DEVICE_ID=1001
MM154 298 60 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3540 $Y=75  $PIN_XY=3570,158,3540,75,3510,158 $DEVICE_ID=1001
MM155 266 59 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3540 $Y=-1072  $PIN_XY=3570,-990,3540,-1072,3510,-990 $DEVICE_ID=1001
MM156 234 58 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3540 $Y=-2219  $PIN_XY=3570,-2136,3540,-2219,3510,-2136 $DEVICE_ID=1001
MM157 18 60 295 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3204 $Y=75  $PIN_XY=3234,158,3204,75,3174,158 $DEVICE_ID=1001
MM158 18 59 263 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3204 $Y=-1072  $PIN_XY=3234,-990,3204,-1072,3174,-990 $DEVICE_ID=1001
MM159 18 58 231 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3204 $Y=-2219  $PIN_XY=3234,-2136,3204,-2219,3174,-2136 $DEVICE_ID=1001
MM160 GND! 296 295 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2868 $Y=304  $PIN_XY=(2898,332,2898,158),2868,304,(2838,332,2838,158) $DEVICE_ID=1001
MM161 GND! 264 263 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2868 $Y=-720  $PIN_XY=(2898,-816,2898,-990),2868,-720,(2838,-816,2838,-990) $DEVICE_ID=1001
MM162 GND! 232 231 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2868 $Y=-1867  $PIN_XY=(2898,-1962,2898,-2136),2868,-1867,(2838,-1962,2838,-2136) $DEVICE_ID=1001
MM163 296 295 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2532 $Y=304  $PIN_XY=(2562,332,2562,158),2532,304,(2502,332,2502,158) $DEVICE_ID=1001
MM164 264 263 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2532 $Y=-720  $PIN_XY=(2562,-816,2562,-990),2532,-720,(2502,-816,2502,-990) $DEVICE_ID=1001
MM165 232 231 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2532 $Y=-1867  $PIN_XY=(2562,-1962,2562,-2136),2532,-1867,(2502,-1962,2502,-2136) $DEVICE_ID=1001
MM166 296 60 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2196 $Y=75  $PIN_XY=2226,158,2196,75,2166,158 $DEVICE_ID=1001
MM167 264 59 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2196 $Y=-1072  $PIN_XY=2226,-990,2196,-1072,2166,-990 $DEVICE_ID=1001
MM168 232 58 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2196 $Y=-2219  $PIN_XY=2226,-2136,2196,-2219,2166,-2136 $DEVICE_ID=1001
MM169 16 60 293 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1860 $Y=75  $PIN_XY=1890,158,1860,75,1830,158 $DEVICE_ID=1001
MM170 16 59 261 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1860 $Y=-1072  $PIN_XY=1890,-990,1860,-1072,1830,-990 $DEVICE_ID=1001
MM171 16 58 229 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1860 $Y=-2219  $PIN_XY=1890,-2136,1860,-2219,1830,-2136 $DEVICE_ID=1001
MM172 GND! 294 293 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1524 $Y=304  $PIN_XY=(1554,332,1554,158),1524,304,(1494,332,1494,158) $DEVICE_ID=1001
MM173 GND! 262 261 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1524 $Y=-720  $PIN_XY=(1554,-816,1554,-990),1524,-720,(1494,-816,1494,-990) $DEVICE_ID=1001
MM174 GND! 230 229 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1524 $Y=-1867  $PIN_XY=(1554,-1962,1554,-2136),1524,-1867,(1494,-1962,1494,-2136) $DEVICE_ID=1001
MM175 294 293 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1188 $Y=304  $PIN_XY=(1218,332,1218,158),1188,304,(1158,332,1158,158) $DEVICE_ID=1001
MM176 262 261 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1188 $Y=-720  $PIN_XY=(1218,-816,1218,-990),1188,-720,(1158,-816,1158,-990) $DEVICE_ID=1001
MM177 230 229 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1188 $Y=-1867  $PIN_XY=(1218,-1962,1218,-2136),1188,-1867,(1158,-1962,1158,-2136) $DEVICE_ID=1001
MM178 294 60 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=852 $Y=75  $PIN_XY=882,158,852,75,822,158 $DEVICE_ID=1001
MM179 262 59 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=852 $Y=-1072  $PIN_XY=882,-990,852,-1072,822,-990 $DEVICE_ID=1001
MM180 230 58 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=852 $Y=-2219  $PIN_XY=882,-2136,852,-2219,822,-2136 $DEVICE_ID=1001
MM181 13 60 291 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=516 $Y=75  $PIN_XY=546,158,516,75,486,158 $DEVICE_ID=1001
MM182 13 59 259 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=516 $Y=-1072  $PIN_XY=546,-990,516,-1072,486,-990 $DEVICE_ID=1001
MM183 13 58 227 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=516 $Y=-2219  $PIN_XY=546,-2136,516,-2219,486,-2136 $DEVICE_ID=1001
MM184 GND! 292 291 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=180 $Y=304  $PIN_XY=(210,332,210,158),180,304,(150,332,150,158) $DEVICE_ID=1001
MM185 GND! 260 259 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=180 $Y=-720  $PIN_XY=(210,-816,210,-990),180,-720,(150,-816,150,-990) $DEVICE_ID=1001
MM186 GND! 228 227 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=180 $Y=-1867  $PIN_XY=(210,-1962,210,-2136),180,-1867,(150,-1962,150,-2136) $DEVICE_ID=1001
MM187 292 291 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=-156 $Y=304  $PIN_XY=(-126,332,-126,158),-156,304,(-186,332,-186,158) $DEVICE_ID=1001
MM188 260 259 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=-156 $Y=-720  $PIN_XY=(-126,-816,-126,-990),-156,-720,(-186,-816,-186,-990) $DEVICE_ID=1001
MM189 228 227 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=-156 $Y=-1867  $PIN_XY=(-126,-1962,-126,-2136),-156,-1867,(-186,-1962,-186,-2136) $DEVICE_ID=1001
MM190 292 60 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=-492 $Y=75  $PIN_XY=-462,158,-492,75,-522,158 $DEVICE_ID=1001
MM191 260 59 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=-492 $Y=-1072  $PIN_XY=-462,-990,-492,-1072,-522,-990 $DEVICE_ID=1001
MM192 228 58 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=-492 $Y=-2219  $PIN_XY=-462,-2136,-492,-2219,-522,-2136 $DEVICE_ID=1001
MM193 44 57 225 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20676 $Y=-3364  $PIN_XY=20706,-3284,20676,-3364,20646,-3284 $DEVICE_ID=1001
MM194 44 56 193 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20676 $Y=-4515  $PIN_XY=20706,-4432,20676,-4515,20646,-4432 $DEVICE_ID=1001
MM195 44 55 161 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20676 $Y=-5662  $PIN_XY=20706,-5580,20676,-5662,20646,-5580 $DEVICE_ID=1001
MM196 GND! 226 225 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=20340 $Y=-3012  $PIN_XY=(20370,-3110,20370,-3284),20340,-3012,(20310,-3110,20310,-3284) $DEVICE_ID=1001
MM197 GND! 194 193 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=20340 $Y=-4160  $PIN_XY=(20370,-4258,20370,-4432),20340,-4160,(20310,-4258,20310,-4432) $DEVICE_ID=1001
MM198 GND! 162 161 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=20340 $Y=-5310  $PIN_XY=(20370,-5406,20370,-5580),20340,-5310,(20310,-5406,20310,-5580) $DEVICE_ID=1001
MM199 226 225 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=20004 $Y=-3012  $PIN_XY=(20034,-3110,20034,-3284),20004,-3012,(19974,-3110,19974,-3284) $DEVICE_ID=1001
MM200 194 193 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=20004 $Y=-4160  $PIN_XY=(20034,-4258,20034,-4432),20004,-4160,(19974,-4258,19974,-4432) $DEVICE_ID=1001
MM201 162 161 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=20004 $Y=-5310  $PIN_XY=(20034,-5406,20034,-5580),20004,-5310,(19974,-5406,19974,-5580) $DEVICE_ID=1001
MM202 226 57 43 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=19668 $Y=-3364  $PIN_XY=19698,-3284,19668,-3364,19638,-3284 $DEVICE_ID=1001
MM203 194 56 43 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=19668 $Y=-4515  $PIN_XY=19698,-4432,19668,-4515,19638,-4432 $DEVICE_ID=1001
MM204 162 55 43 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=19668 $Y=-5662  $PIN_XY=19698,-5580,19668,-5662,19638,-5580 $DEVICE_ID=1001
MM205 42 57 223 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=19332 $Y=-3364  $PIN_XY=19362,-3284,19332,-3364,19302,-3284 $DEVICE_ID=1001
MM206 42 56 191 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=19332 $Y=-4515  $PIN_XY=19362,-4432,19332,-4515,19302,-4432 $DEVICE_ID=1001
MM207 42 55 159 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=19332 $Y=-5662  $PIN_XY=19362,-5580,19332,-5662,19302,-5580 $DEVICE_ID=1001
MM208 GND! 224 223 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=18996 $Y=-3012  $PIN_XY=(19026,-3110,19026,-3284),18996,-3012,(18966,-3110,18966,-3284) $DEVICE_ID=1001
MM209 GND! 192 191 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=18996 $Y=-4160  $PIN_XY=(19026,-4258,19026,-4432),18996,-4160,(18966,-4258,18966,-4432) $DEVICE_ID=1001
MM210 GND! 160 159 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=18996 $Y=-5310  $PIN_XY=(19026,-5406,19026,-5580),18996,-5310,(18966,-5406,18966,-5580) $DEVICE_ID=1001
MM211 224 223 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=18660 $Y=-3012  $PIN_XY=(18690,-3110,18690,-3284),18660,-3012,(18630,-3110,18630,-3284) $DEVICE_ID=1001
MM212 192 191 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=18660 $Y=-4160  $PIN_XY=(18690,-4258,18690,-4432),18660,-4160,(18630,-4258,18630,-4432) $DEVICE_ID=1001
MM213 160 159 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=18660 $Y=-5310  $PIN_XY=(18690,-5406,18690,-5580),18660,-5310,(18630,-5406,18630,-5580) $DEVICE_ID=1001
MM214 224 57 41 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18324 $Y=-3364  $PIN_XY=18354,-3284,18324,-3364,18294,-3284 $DEVICE_ID=1001
MM215 192 56 41 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18324 $Y=-4515  $PIN_XY=18354,-4432,18324,-4515,18294,-4432 $DEVICE_ID=1001
MM216 160 55 41 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18324 $Y=-5662  $PIN_XY=18354,-5580,18324,-5662,18294,-5580 $DEVICE_ID=1001
MM217 40 57 221 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17988 $Y=-3364  $PIN_XY=18018,-3284,17988,-3364,17958,-3284 $DEVICE_ID=1001
MM218 40 56 189 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17988 $Y=-4515  $PIN_XY=18018,-4432,17988,-4515,17958,-4432 $DEVICE_ID=1001
MM219 40 55 157 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17988 $Y=-5662  $PIN_XY=18018,-5580,17988,-5662,17958,-5580 $DEVICE_ID=1001
MM220 GND! 222 221 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17652 $Y=-3012  $PIN_XY=(17682,-3110,17682,-3284),17652,-3012,(17622,-3110,17622,-3284) $DEVICE_ID=1001
MM221 GND! 190 189 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17652 $Y=-4160  $PIN_XY=(17682,-4258,17682,-4432),17652,-4160,(17622,-4258,17622,-4432) $DEVICE_ID=1001
MM222 GND! 158 157 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17652 $Y=-5310  $PIN_XY=(17682,-5406,17682,-5580),17652,-5310,(17622,-5406,17622,-5580) $DEVICE_ID=1001
MM223 222 221 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17316 $Y=-3012  $PIN_XY=(17346,-3110,17346,-3284),17316,-3012,(17286,-3110,17286,-3284) $DEVICE_ID=1001
MM224 190 189 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17316 $Y=-4160  $PIN_XY=(17346,-4258,17346,-4432),17316,-4160,(17286,-4258,17286,-4432) $DEVICE_ID=1001
MM225 158 157 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17316 $Y=-5310  $PIN_XY=(17346,-5406,17346,-5580),17316,-5310,(17286,-5406,17286,-5580) $DEVICE_ID=1001
MM226 222 57 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16980 $Y=-3364  $PIN_XY=17010,-3284,16980,-3364,16950,-3284 $DEVICE_ID=1001
MM227 190 56 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16980 $Y=-4515  $PIN_XY=17010,-4432,16980,-4515,16950,-4432 $DEVICE_ID=1001
MM228 158 55 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16980 $Y=-5662  $PIN_XY=17010,-5580,16980,-5662,16950,-5580 $DEVICE_ID=1001
MM229 38 57 219 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16644 $Y=-3364  $PIN_XY=16674,-3284,16644,-3364,16614,-3284 $DEVICE_ID=1001
MM230 38 56 187 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16644 $Y=-4515  $PIN_XY=16674,-4432,16644,-4515,16614,-4432 $DEVICE_ID=1001
MM231 38 55 155 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16644 $Y=-5662  $PIN_XY=16674,-5580,16644,-5662,16614,-5580 $DEVICE_ID=1001
MM232 GND! 220 219 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=16308 $Y=-3012  $PIN_XY=(16338,-3110,16338,-3284),16308,-3012,(16278,-3110,16278,-3284) $DEVICE_ID=1001
MM233 GND! 188 187 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=16308 $Y=-4160  $PIN_XY=(16338,-4258,16338,-4432),16308,-4160,(16278,-4258,16278,-4432) $DEVICE_ID=1001
MM234 GND! 156 155 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=16308 $Y=-5310  $PIN_XY=(16338,-5406,16338,-5580),16308,-5310,(16278,-5406,16278,-5580) $DEVICE_ID=1001
MM235 220 219 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=15972 $Y=-3012  $PIN_XY=(16002,-3110,16002,-3284),15972,-3012,(15942,-3110,15942,-3284) $DEVICE_ID=1001
MM236 188 187 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=15972 $Y=-4160  $PIN_XY=(16002,-4258,16002,-4432),15972,-4160,(15942,-4258,15942,-4432) $DEVICE_ID=1001
MM237 156 155 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=15972 $Y=-5310  $PIN_XY=(16002,-5406,16002,-5580),15972,-5310,(15942,-5406,15942,-5580) $DEVICE_ID=1001
MM238 220 57 37 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15636 $Y=-3364  $PIN_XY=15666,-3284,15636,-3364,15606,-3284 $DEVICE_ID=1001
MM239 188 56 37 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15636 $Y=-4515  $PIN_XY=15666,-4432,15636,-4515,15606,-4432 $DEVICE_ID=1001
MM240 156 55 37 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15636 $Y=-5662  $PIN_XY=15666,-5580,15636,-5662,15606,-5580 $DEVICE_ID=1001
MM241 36 57 217 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15300 $Y=-3364  $PIN_XY=15330,-3284,15300,-3364,15270,-3284 $DEVICE_ID=1001
MM242 36 56 185 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15300 $Y=-4515  $PIN_XY=15330,-4432,15300,-4515,15270,-4432 $DEVICE_ID=1001
MM243 36 55 153 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15300 $Y=-5662  $PIN_XY=15330,-5580,15300,-5662,15270,-5580 $DEVICE_ID=1001
MM244 GND! 218 217 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14964 $Y=-3012  $PIN_XY=(14994,-3110,14994,-3284),14964,-3012,(14934,-3110,14934,-3284) $DEVICE_ID=1001
MM245 GND! 186 185 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14964 $Y=-4160  $PIN_XY=(14994,-4258,14994,-4432),14964,-4160,(14934,-4258,14934,-4432) $DEVICE_ID=1001
MM246 GND! 154 153 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14964 $Y=-5310  $PIN_XY=(14994,-5406,14994,-5580),14964,-5310,(14934,-5406,14934,-5580) $DEVICE_ID=1001
MM247 218 217 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14628 $Y=-3012  $PIN_XY=(14658,-3110,14658,-3284),14628,-3012,(14598,-3110,14598,-3284) $DEVICE_ID=1001
MM248 186 185 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14628 $Y=-4160  $PIN_XY=(14658,-4258,14658,-4432),14628,-4160,(14598,-4258,14598,-4432) $DEVICE_ID=1001
MM249 154 153 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14628 $Y=-5310  $PIN_XY=(14658,-5406,14658,-5580),14628,-5310,(14598,-5406,14598,-5580) $DEVICE_ID=1001
MM250 218 57 35 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14292 $Y=-3364  $PIN_XY=14322,-3284,14292,-3364,14262,-3284 $DEVICE_ID=1001
MM251 186 56 35 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14292 $Y=-4515  $PIN_XY=14322,-4432,14292,-4515,14262,-4432 $DEVICE_ID=1001
MM252 154 55 35 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14292 $Y=-5662  $PIN_XY=14322,-5580,14292,-5662,14262,-5580 $DEVICE_ID=1001
MM253 34 57 215 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13956 $Y=-3364  $PIN_XY=13986,-3284,13956,-3364,13926,-3284 $DEVICE_ID=1001
MM254 34 56 183 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13956 $Y=-4515  $PIN_XY=13986,-4432,13956,-4515,13926,-4432 $DEVICE_ID=1001
MM255 34 55 151 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13956 $Y=-5662  $PIN_XY=13986,-5580,13956,-5662,13926,-5580 $DEVICE_ID=1001
MM256 GND! 216 215 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13620 $Y=-3012  $PIN_XY=(13650,-3110,13650,-3284),13620,-3012,(13590,-3110,13590,-3284) $DEVICE_ID=1001
MM257 GND! 184 183 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13620 $Y=-4160  $PIN_XY=(13650,-4258,13650,-4432),13620,-4160,(13590,-4258,13590,-4432) $DEVICE_ID=1001
MM258 GND! 152 151 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13620 $Y=-5310  $PIN_XY=(13650,-5406,13650,-5580),13620,-5310,(13590,-5406,13590,-5580) $DEVICE_ID=1001
MM259 216 215 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13284 $Y=-3012  $PIN_XY=(13314,-3110,13314,-3284),13284,-3012,(13254,-3110,13254,-3284) $DEVICE_ID=1001
MM260 184 183 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13284 $Y=-4160  $PIN_XY=(13314,-4258,13314,-4432),13284,-4160,(13254,-4258,13254,-4432) $DEVICE_ID=1001
MM261 152 151 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13284 $Y=-5310  $PIN_XY=(13314,-5406,13314,-5580),13284,-5310,(13254,-5406,13254,-5580) $DEVICE_ID=1001
MM262 216 57 33 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12948 $Y=-3364  $PIN_XY=12978,-3284,12948,-3364,12918,-3284 $DEVICE_ID=1001
MM263 184 56 33 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12948 $Y=-4515  $PIN_XY=12978,-4432,12948,-4515,12918,-4432 $DEVICE_ID=1001
MM264 152 55 33 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12948 $Y=-5662  $PIN_XY=12978,-5580,12948,-5662,12918,-5580 $DEVICE_ID=1001
MM265 32 57 213 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12612 $Y=-3364  $PIN_XY=12642,-3284,12612,-3364,12582,-3284 $DEVICE_ID=1001
MM266 32 56 181 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12612 $Y=-4515  $PIN_XY=12642,-4432,12612,-4515,12582,-4432 $DEVICE_ID=1001
MM267 32 55 149 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12612 $Y=-5662  $PIN_XY=12642,-5580,12612,-5662,12582,-5580 $DEVICE_ID=1001
MM268 GND! 214 213 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=12276 $Y=-3012  $PIN_XY=(12306,-3110,12306,-3284),12276,-3012,(12246,-3110,12246,-3284) $DEVICE_ID=1001
MM269 GND! 182 181 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=12276 $Y=-4160  $PIN_XY=(12306,-4258,12306,-4432),12276,-4160,(12246,-4258,12246,-4432) $DEVICE_ID=1001
MM270 GND! 150 149 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=12276 $Y=-5310  $PIN_XY=(12306,-5406,12306,-5580),12276,-5310,(12246,-5406,12246,-5580) $DEVICE_ID=1001
MM271 214 213 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11940 $Y=-3012  $PIN_XY=(11970,-3110,11970,-3284),11940,-3012,(11910,-3110,11910,-3284) $DEVICE_ID=1001
MM272 182 181 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11940 $Y=-4160  $PIN_XY=(11970,-4258,11970,-4432),11940,-4160,(11910,-4258,11910,-4432) $DEVICE_ID=1001
MM273 150 149 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11940 $Y=-5310  $PIN_XY=(11970,-5406,11970,-5580),11940,-5310,(11910,-5406,11910,-5580) $DEVICE_ID=1001
MM274 214 57 31 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11604 $Y=-3364  $PIN_XY=11634,-3284,11604,-3364,11574,-3284 $DEVICE_ID=1001
MM275 182 56 31 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11604 $Y=-4515  $PIN_XY=11634,-4432,11604,-4515,11574,-4432 $DEVICE_ID=1001
MM276 150 55 31 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11604 $Y=-5662  $PIN_XY=11634,-5580,11604,-5662,11574,-5580 $DEVICE_ID=1001
MM277 30 57 211 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11268 $Y=-3364  $PIN_XY=11298,-3284,11268,-3364,11238,-3284 $DEVICE_ID=1001
MM278 30 56 179 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11268 $Y=-4515  $PIN_XY=11298,-4432,11268,-4515,11238,-4432 $DEVICE_ID=1001
MM279 30 55 147 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11268 $Y=-5662  $PIN_XY=11298,-5580,11268,-5662,11238,-5580 $DEVICE_ID=1001
MM280 GND! 212 211 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10932 $Y=-3012  $PIN_XY=(10962,-3110,10962,-3284),10932,-3012,(10902,-3110,10902,-3284) $DEVICE_ID=1001
MM281 GND! 180 179 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10932 $Y=-4160  $PIN_XY=(10962,-4258,10962,-4432),10932,-4160,(10902,-4258,10902,-4432) $DEVICE_ID=1001
MM282 GND! 148 147 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10932 $Y=-5310  $PIN_XY=(10962,-5406,10962,-5580),10932,-5310,(10902,-5406,10902,-5580) $DEVICE_ID=1001
MM283 212 211 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10596 $Y=-3012  $PIN_XY=(10626,-3110,10626,-3284),10596,-3012,(10566,-3110,10566,-3284) $DEVICE_ID=1001
MM284 180 179 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10596 $Y=-4160  $PIN_XY=(10626,-4258,10626,-4432),10596,-4160,(10566,-4258,10566,-4432) $DEVICE_ID=1001
MM285 148 147 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10596 $Y=-5310  $PIN_XY=(10626,-5406,10626,-5580),10596,-5310,(10566,-5406,10566,-5580) $DEVICE_ID=1001
MM286 212 57 29 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10260 $Y=-3364  $PIN_XY=10290,-3284,10260,-3364,10230,-3284 $DEVICE_ID=1001
MM287 180 56 29 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10260 $Y=-4515  $PIN_XY=10290,-4432,10260,-4515,10230,-4432 $DEVICE_ID=1001
MM288 148 55 29 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10260 $Y=-5662  $PIN_XY=10290,-5580,10260,-5662,10230,-5580 $DEVICE_ID=1001
MM289 28 57 209 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9924 $Y=-3364  $PIN_XY=9954,-3284,9924,-3364,9894,-3284 $DEVICE_ID=1001
MM290 28 56 177 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9924 $Y=-4515  $PIN_XY=9954,-4432,9924,-4515,9894,-4432 $DEVICE_ID=1001
MM291 28 55 145 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9924 $Y=-5662  $PIN_XY=9954,-5580,9924,-5662,9894,-5580 $DEVICE_ID=1001
MM292 GND! 210 209 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9588 $Y=-3012  $PIN_XY=(9618,-3110,9618,-3284),9588,-3012,(9558,-3110,9558,-3284) $DEVICE_ID=1001
MM293 GND! 178 177 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9588 $Y=-4160  $PIN_XY=(9618,-4258,9618,-4432),9588,-4160,(9558,-4258,9558,-4432) $DEVICE_ID=1001
MM294 GND! 146 145 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9588 $Y=-5310  $PIN_XY=(9618,-5406,9618,-5580),9588,-5310,(9558,-5406,9558,-5580) $DEVICE_ID=1001
MM295 210 209 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9252 $Y=-3012  $PIN_XY=(9282,-3110,9282,-3284),9252,-3012,(9222,-3110,9222,-3284) $DEVICE_ID=1001
MM296 178 177 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9252 $Y=-4160  $PIN_XY=(9282,-4258,9282,-4432),9252,-4160,(9222,-4258,9222,-4432) $DEVICE_ID=1001
MM297 146 145 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9252 $Y=-5310  $PIN_XY=(9282,-5406,9282,-5580),9252,-5310,(9222,-5406,9222,-5580) $DEVICE_ID=1001
MM298 210 57 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8916 $Y=-3364  $PIN_XY=8946,-3284,8916,-3364,8886,-3284 $DEVICE_ID=1001
MM299 178 56 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8916 $Y=-4515  $PIN_XY=8946,-4432,8916,-4515,8886,-4432 $DEVICE_ID=1001
MM300 146 55 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8916 $Y=-5662  $PIN_XY=8946,-5580,8916,-5662,8886,-5580 $DEVICE_ID=1001
MM301 26 57 207 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8580 $Y=-3364  $PIN_XY=8610,-3284,8580,-3364,8550,-3284 $DEVICE_ID=1001
MM302 26 56 175 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8580 $Y=-4515  $PIN_XY=8610,-4432,8580,-4515,8550,-4432 $DEVICE_ID=1001
MM303 26 55 143 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8580 $Y=-5662  $PIN_XY=8610,-5580,8580,-5662,8550,-5580 $DEVICE_ID=1001
MM304 GND! 208 207 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8244 $Y=-3012  $PIN_XY=(8274,-3110,8274,-3284),8244,-3012,(8214,-3110,8214,-3284) $DEVICE_ID=1001
MM305 GND! 176 175 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8244 $Y=-4160  $PIN_XY=(8274,-4258,8274,-4432),8244,-4160,(8214,-4258,8214,-4432) $DEVICE_ID=1001
MM306 GND! 144 143 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8244 $Y=-5310  $PIN_XY=(8274,-5406,8274,-5580),8244,-5310,(8214,-5406,8214,-5580) $DEVICE_ID=1001
MM307 208 207 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7908 $Y=-3012  $PIN_XY=(7938,-3110,7938,-3284),7908,-3012,(7878,-3110,7878,-3284) $DEVICE_ID=1001
MM308 176 175 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7908 $Y=-4160  $PIN_XY=(7938,-4258,7938,-4432),7908,-4160,(7878,-4258,7878,-4432) $DEVICE_ID=1001
MM309 144 143 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7908 $Y=-5310  $PIN_XY=(7938,-5406,7938,-5580),7908,-5310,(7878,-5406,7878,-5580) $DEVICE_ID=1001
MM310 208 57 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7572 $Y=-3364  $PIN_XY=7602,-3284,7572,-3364,7542,-3284 $DEVICE_ID=1001
MM311 176 56 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7572 $Y=-4515  $PIN_XY=7602,-4432,7572,-4515,7542,-4432 $DEVICE_ID=1001
MM312 144 55 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7572 $Y=-5662  $PIN_XY=7602,-5580,7572,-5662,7542,-5580 $DEVICE_ID=1001
MM313 24 57 205 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7236 $Y=-3364  $PIN_XY=7266,-3284,7236,-3364,7206,-3284 $DEVICE_ID=1001
MM314 24 56 173 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7236 $Y=-4515  $PIN_XY=7266,-4432,7236,-4515,7206,-4432 $DEVICE_ID=1001
MM315 24 55 141 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7236 $Y=-5662  $PIN_XY=7266,-5580,7236,-5662,7206,-5580 $DEVICE_ID=1001
MM316 GND! 206 205 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6900 $Y=-3012  $PIN_XY=(6930,-3110,6930,-3284),6900,-3012,(6870,-3110,6870,-3284) $DEVICE_ID=1001
MM317 GND! 174 173 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6900 $Y=-4160  $PIN_XY=(6930,-4258,6930,-4432),6900,-4160,(6870,-4258,6870,-4432) $DEVICE_ID=1001
MM318 GND! 142 141 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6900 $Y=-5310  $PIN_XY=(6930,-5406,6930,-5580),6900,-5310,(6870,-5406,6870,-5580) $DEVICE_ID=1001
MM319 206 205 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6564 $Y=-3012  $PIN_XY=(6594,-3110,6594,-3284),6564,-3012,(6534,-3110,6534,-3284) $DEVICE_ID=1001
MM320 174 173 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6564 $Y=-4160  $PIN_XY=(6594,-4258,6594,-4432),6564,-4160,(6534,-4258,6534,-4432) $DEVICE_ID=1001
MM321 142 141 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6564 $Y=-5310  $PIN_XY=(6594,-5406,6594,-5580),6564,-5310,(6534,-5406,6534,-5580) $DEVICE_ID=1001
MM322 206 57 23 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6228 $Y=-3364  $PIN_XY=6258,-3284,6228,-3364,6198,-3284 $DEVICE_ID=1001
MM323 174 56 23 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6228 $Y=-4515  $PIN_XY=6258,-4432,6228,-4515,6198,-4432 $DEVICE_ID=1001
MM324 142 55 23 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6228 $Y=-5662  $PIN_XY=6258,-5580,6228,-5662,6198,-5580 $DEVICE_ID=1001
MM325 22 57 203 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5892 $Y=-3364  $PIN_XY=5922,-3284,5892,-3364,5862,-3284 $DEVICE_ID=1001
MM326 22 56 171 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5892 $Y=-4515  $PIN_XY=5922,-4432,5892,-4515,5862,-4432 $DEVICE_ID=1001
MM327 22 55 139 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5892 $Y=-5662  $PIN_XY=5922,-5580,5892,-5662,5862,-5580 $DEVICE_ID=1001
MM328 GND! 204 203 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5556 $Y=-3012  $PIN_XY=(5586,-3110,5586,-3284),5556,-3012,(5526,-3110,5526,-3284) $DEVICE_ID=1001
MM329 GND! 172 171 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5556 $Y=-4160  $PIN_XY=(5586,-4258,5586,-4432),5556,-4160,(5526,-4258,5526,-4432) $DEVICE_ID=1001
MM330 GND! 140 139 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5556 $Y=-5310  $PIN_XY=(5586,-5406,5586,-5580),5556,-5310,(5526,-5406,5526,-5580) $DEVICE_ID=1001
MM331 204 203 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5220 $Y=-3012  $PIN_XY=(5250,-3110,5250,-3284),5220,-3012,(5190,-3110,5190,-3284) $DEVICE_ID=1001
MM332 172 171 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5220 $Y=-4160  $PIN_XY=(5250,-4258,5250,-4432),5220,-4160,(5190,-4258,5190,-4432) $DEVICE_ID=1001
MM333 140 139 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5220 $Y=-5310  $PIN_XY=(5250,-5406,5250,-5580),5220,-5310,(5190,-5406,5190,-5580) $DEVICE_ID=1001
MM334 204 57 21 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4884 $Y=-3364  $PIN_XY=4914,-3284,4884,-3364,4854,-3284 $DEVICE_ID=1001
MM335 172 56 21 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4884 $Y=-4515  $PIN_XY=4914,-4432,4884,-4515,4854,-4432 $DEVICE_ID=1001
MM336 140 55 21 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4884 $Y=-5662  $PIN_XY=4914,-5580,4884,-5662,4854,-5580 $DEVICE_ID=1001
MM337 20 57 201 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4548 $Y=-3364  $PIN_XY=4578,-3284,4548,-3364,4518,-3284 $DEVICE_ID=1001
MM338 20 56 169 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4548 $Y=-4515  $PIN_XY=4578,-4432,4548,-4515,4518,-4432 $DEVICE_ID=1001
MM339 20 55 137 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4548 $Y=-5662  $PIN_XY=4578,-5580,4548,-5662,4518,-5580 $DEVICE_ID=1001
MM340 GND! 202 201 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4212 $Y=-3012  $PIN_XY=(4242,-3110,4242,-3284),4212,-3012,(4182,-3110,4182,-3284) $DEVICE_ID=1001
MM341 GND! 170 169 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4212 $Y=-4160  $PIN_XY=(4242,-4258,4242,-4432),4212,-4160,(4182,-4258,4182,-4432) $DEVICE_ID=1001
MM342 GND! 138 137 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4212 $Y=-5310  $PIN_XY=(4242,-5406,4242,-5580),4212,-5310,(4182,-5406,4182,-5580) $DEVICE_ID=1001
MM343 202 201 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3876 $Y=-3012  $PIN_XY=(3906,-3110,3906,-3284),3876,-3012,(3846,-3110,3846,-3284) $DEVICE_ID=1001
MM344 170 169 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3876 $Y=-4160  $PIN_XY=(3906,-4258,3906,-4432),3876,-4160,(3846,-4258,3846,-4432) $DEVICE_ID=1001
MM345 138 137 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3876 $Y=-5310  $PIN_XY=(3906,-5406,3906,-5580),3876,-5310,(3846,-5406,3846,-5580) $DEVICE_ID=1001
MM346 202 57 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3540 $Y=-3364  $PIN_XY=3570,-3284,3540,-3364,3510,-3284 $DEVICE_ID=1001
MM347 170 56 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3540 $Y=-4515  $PIN_XY=3570,-4432,3540,-4515,3510,-4432 $DEVICE_ID=1001
MM348 138 55 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3540 $Y=-5662  $PIN_XY=3570,-5580,3540,-5662,3510,-5580 $DEVICE_ID=1001
MM349 18 57 199 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3204 $Y=-3364  $PIN_XY=3234,-3284,3204,-3364,3174,-3284 $DEVICE_ID=1001
MM350 18 56 167 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3204 $Y=-4515  $PIN_XY=3234,-4432,3204,-4515,3174,-4432 $DEVICE_ID=1001
MM351 18 55 135 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3204 $Y=-5662  $PIN_XY=3234,-5580,3204,-5662,3174,-5580 $DEVICE_ID=1001
MM352 GND! 200 199 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2868 $Y=-3012  $PIN_XY=(2898,-3110,2898,-3284),2868,-3012,(2838,-3110,2838,-3284) $DEVICE_ID=1001
MM353 GND! 168 167 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2868 $Y=-4160  $PIN_XY=(2898,-4258,2898,-4432),2868,-4160,(2838,-4258,2838,-4432) $DEVICE_ID=1001
MM354 GND! 136 135 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2868 $Y=-5310  $PIN_XY=(2898,-5406,2898,-5580),2868,-5310,(2838,-5406,2838,-5580) $DEVICE_ID=1001
MM355 200 199 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2532 $Y=-3012  $PIN_XY=(2562,-3110,2562,-3284),2532,-3012,(2502,-3110,2502,-3284) $DEVICE_ID=1001
MM356 168 167 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2532 $Y=-4160  $PIN_XY=(2562,-4258,2562,-4432),2532,-4160,(2502,-4258,2502,-4432) $DEVICE_ID=1001
MM357 136 135 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2532 $Y=-5310  $PIN_XY=(2562,-5406,2562,-5580),2532,-5310,(2502,-5406,2502,-5580) $DEVICE_ID=1001
MM358 200 57 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2196 $Y=-3364  $PIN_XY=2226,-3284,2196,-3364,2166,-3284 $DEVICE_ID=1001
MM359 168 56 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2196 $Y=-4515  $PIN_XY=2226,-4432,2196,-4515,2166,-4432 $DEVICE_ID=1001
MM360 136 55 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2196 $Y=-5662  $PIN_XY=2226,-5580,2196,-5662,2166,-5580 $DEVICE_ID=1001
MM361 16 57 197 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1860 $Y=-3364  $PIN_XY=1890,-3284,1860,-3364,1830,-3284 $DEVICE_ID=1001
MM362 16 56 165 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1860 $Y=-4515  $PIN_XY=1890,-4432,1860,-4515,1830,-4432 $DEVICE_ID=1001
MM363 16 55 133 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1860 $Y=-5662  $PIN_XY=1890,-5580,1860,-5662,1830,-5580 $DEVICE_ID=1001
MM364 GND! 198 197 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1524 $Y=-3012  $PIN_XY=(1554,-3110,1554,-3284),1524,-3012,(1494,-3110,1494,-3284) $DEVICE_ID=1001
MM365 GND! 166 165 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1524 $Y=-4160  $PIN_XY=(1554,-4258,1554,-4432),1524,-4160,(1494,-4258,1494,-4432) $DEVICE_ID=1001
MM366 GND! 134 133 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1524 $Y=-5310  $PIN_XY=(1554,-5406,1554,-5580),1524,-5310,(1494,-5406,1494,-5580) $DEVICE_ID=1001
MM367 198 197 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1188 $Y=-3012  $PIN_XY=(1218,-3110,1218,-3284),1188,-3012,(1158,-3110,1158,-3284) $DEVICE_ID=1001
MM368 166 165 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1188 $Y=-4160  $PIN_XY=(1218,-4258,1218,-4432),1188,-4160,(1158,-4258,1158,-4432) $DEVICE_ID=1001
MM369 134 133 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1188 $Y=-5310  $PIN_XY=(1218,-5406,1218,-5580),1188,-5310,(1158,-5406,1158,-5580) $DEVICE_ID=1001
MM370 198 57 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=852 $Y=-3364  $PIN_XY=882,-3284,852,-3364,822,-3284 $DEVICE_ID=1001
MM371 166 56 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=852 $Y=-4515  $PIN_XY=882,-4432,852,-4515,822,-4432 $DEVICE_ID=1001
MM372 134 55 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=852 $Y=-5662  $PIN_XY=882,-5580,852,-5662,822,-5580 $DEVICE_ID=1001
MM373 13 57 195 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=516 $Y=-3364  $PIN_XY=546,-3284,516,-3364,486,-3284 $DEVICE_ID=1001
MM374 13 56 163 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=516 $Y=-4515  $PIN_XY=546,-4432,516,-4515,486,-4432 $DEVICE_ID=1001
MM375 13 55 131 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=516 $Y=-5662  $PIN_XY=546,-5580,516,-5662,486,-5580 $DEVICE_ID=1001
MM376 GND! 196 195 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=180 $Y=-3012  $PIN_XY=(210,-3110,210,-3284),180,-3012,(150,-3110,150,-3284) $DEVICE_ID=1001
MM377 GND! 164 163 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=180 $Y=-4160  $PIN_XY=(210,-4258,210,-4432),180,-4160,(150,-4258,150,-4432) $DEVICE_ID=1001
MM378 GND! 132 131 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=180 $Y=-5310  $PIN_XY=(210,-5406,210,-5580),180,-5310,(150,-5406,150,-5580) $DEVICE_ID=1001
MM379 196 195 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=-156 $Y=-3012  $PIN_XY=(-126,-3110,-126,-3284),-156,-3012,(-186,-3110,-186,-3284) $DEVICE_ID=1001
MM380 164 163 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=-156 $Y=-4160  $PIN_XY=(-126,-4258,-126,-4432),-156,-4160,(-186,-4258,-186,-4432) $DEVICE_ID=1001
MM381 132 131 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=-156 $Y=-5310  $PIN_XY=(-126,-5406,-126,-5580),-156,-5310,(-186,-5406,-186,-5580) $DEVICE_ID=1001
MM382 196 57 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=-492 $Y=-3364  $PIN_XY=-462,-3284,-492,-3364,-522,-3284 $DEVICE_ID=1001
MM383 164 56 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=-492 $Y=-4515  $PIN_XY=-462,-4432,-492,-4515,-522,-4432 $DEVICE_ID=1001
MM384 132 55 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=-492 $Y=-5662  $PIN_XY=-462,-5580,-492,-5662,-522,-5580 $DEVICE_ID=1001
MM385 44 54 129 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20676 $Y=-6809  $PIN_XY=20706,-6726,20676,-6809,20646,-6726 $DEVICE_ID=1001
MM386 44 53 97 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20676 $Y=-7933  $PIN_XY=20706,-7874,20676,-7933,20646,-7874 $DEVICE_ID=1001
MM387 GND! 130 129 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=20340 $Y=-6457  $PIN_XY=(20370,-6552,20370,-6726),20340,-6457,(20310,-6552,20310,-6726) $DEVICE_ID=1001
MM388 GND! 98 97 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=20340 $Y=-7581  $PIN_XY=(20370,-7700,20370,-7874),20340,-7581,(20310,-7700,20310,-7874) $DEVICE_ID=1001
MM389 130 129 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=20004 $Y=-6457  $PIN_XY=(20034,-6552,20034,-6726),20004,-6457,(19974,-6552,19974,-6726) $DEVICE_ID=1001
MM390 98 97 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=20004 $Y=-7581  $PIN_XY=(20034,-7700,20034,-7874),20004,-7581,(19974,-7700,19974,-7874) $DEVICE_ID=1001
MM391 130 54 43 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=19668 $Y=-6809  $PIN_XY=19698,-6726,19668,-6809,19638,-6726 $DEVICE_ID=1001
MM392 98 53 43 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=19668 $Y=-7933  $PIN_XY=19698,-7874,19668,-7933,19638,-7874 $DEVICE_ID=1001
MM393 42 54 127 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=19332 $Y=-6809  $PIN_XY=19362,-6726,19332,-6809,19302,-6726 $DEVICE_ID=1001
MM394 42 53 95 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=19332 $Y=-7933  $PIN_XY=19362,-7874,19332,-7933,19302,-7874 $DEVICE_ID=1001
MM395 GND! 128 127 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=18996 $Y=-6457  $PIN_XY=(19026,-6552,19026,-6726),18996,-6457,(18966,-6552,18966,-6726) $DEVICE_ID=1001
MM396 GND! 96 95 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=18996 $Y=-7596  $PIN_XY=(19026,-7700,19026,-7874),18996,-7596,(18966,-7700,18966,-7874) $DEVICE_ID=1001
MM397 128 127 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=18660 $Y=-6457  $PIN_XY=(18690,-6552,18690,-6726),18660,-6457,(18630,-6552,18630,-6726) $DEVICE_ID=1001
MM398 96 95 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=18660 $Y=-7581  $PIN_XY=(18690,-7700,18690,-7874),18660,-7581,(18630,-7700,18630,-7874) $DEVICE_ID=1001
MM399 128 54 41 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18324 $Y=-6809  $PIN_XY=18354,-6726,18324,-6809,18294,-6726 $DEVICE_ID=1001
MM400 96 53 41 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18324 $Y=-7933  $PIN_XY=18354,-7874,18324,-7933,18294,-7874 $DEVICE_ID=1001
MM401 40 54 125 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17988 $Y=-6809  $PIN_XY=18018,-6726,17988,-6809,17958,-6726 $DEVICE_ID=1001
MM402 40 53 93 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17988 $Y=-7933  $PIN_XY=18018,-7874,17988,-7933,17958,-7874 $DEVICE_ID=1001
MM403 GND! 126 125 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17652 $Y=-6457  $PIN_XY=(17682,-6552,17682,-6726),17652,-6457,(17622,-6552,17622,-6726) $DEVICE_ID=1001
MM404 GND! 94 93 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17652 $Y=-7581  $PIN_XY=(17682,-7700,17682,-7874),17652,-7581,(17622,-7700,17622,-7874) $DEVICE_ID=1001
MM405 126 125 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17316 $Y=-6457  $PIN_XY=(17346,-6552,17346,-6726),17316,-6457,(17286,-6552,17286,-6726) $DEVICE_ID=1001
MM406 94 93 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=17316 $Y=-7581  $PIN_XY=(17346,-7700,17346,-7874),17316,-7581,(17286,-7700,17286,-7874) $DEVICE_ID=1001
MM407 126 54 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16980 $Y=-6809  $PIN_XY=17010,-6726,16980,-6809,16950,-6726 $DEVICE_ID=1001
MM408 94 53 39 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16980 $Y=-7933  $PIN_XY=17010,-7874,16980,-7933,16950,-7874 $DEVICE_ID=1001
MM409 38 54 123 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16644 $Y=-6809  $PIN_XY=16674,-6726,16644,-6809,16614,-6726 $DEVICE_ID=1001
MM410 38 53 91 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16644 $Y=-7933  $PIN_XY=16674,-7874,16644,-7933,16614,-7874 $DEVICE_ID=1001
MM411 GND! 124 123 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=16308 $Y=-6457  $PIN_XY=(16338,-6552,16338,-6726),16308,-6457,(16278,-6552,16278,-6726) $DEVICE_ID=1001
MM412 GND! 92 91 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=16308 $Y=-7581  $PIN_XY=(16338,-7700,16338,-7874),16308,-7581,(16278,-7700,16278,-7874) $DEVICE_ID=1001
MM413 124 123 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=15972 $Y=-6457  $PIN_XY=(16002,-6552,16002,-6726),15972,-6457,(15942,-6552,15942,-6726) $DEVICE_ID=1001
MM414 92 91 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=15972 $Y=-7581  $PIN_XY=(16002,-7700,16002,-7874),15972,-7581,(15942,-7700,15942,-7874) $DEVICE_ID=1001
MM415 124 54 37 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15636 $Y=-6809  $PIN_XY=15666,-6726,15636,-6809,15606,-6726 $DEVICE_ID=1001
MM416 92 53 37 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15636 $Y=-7933  $PIN_XY=15666,-7874,15636,-7933,15606,-7874 $DEVICE_ID=1001
MM417 36 54 121 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15300 $Y=-6809  $PIN_XY=15330,-6726,15300,-6809,15270,-6726 $DEVICE_ID=1001
MM418 36 53 89 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15300 $Y=-7933  $PIN_XY=15330,-7874,15300,-7933,15270,-7874 $DEVICE_ID=1001
MM419 GND! 122 121 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14964 $Y=-6457  $PIN_XY=(14994,-6552,14994,-6726),14964,-6457,(14934,-6552,14934,-6726) $DEVICE_ID=1001
MM420 GND! 90 89 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14964 $Y=-7581  $PIN_XY=(14994,-7700,14994,-7874),14964,-7581,(14934,-7700,14934,-7874) $DEVICE_ID=1001
MM421 122 121 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14628 $Y=-6457  $PIN_XY=(14658,-6552,14658,-6726),14628,-6457,(14598,-6552,14598,-6726) $DEVICE_ID=1001
MM422 90 89 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=14628 $Y=-7581  $PIN_XY=(14658,-7700,14658,-7874),14628,-7581,(14598,-7700,14598,-7874) $DEVICE_ID=1001
MM423 122 54 35 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14292 $Y=-6809  $PIN_XY=14322,-6726,14292,-6809,14262,-6726 $DEVICE_ID=1001
MM424 90 53 35 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14292 $Y=-7933  $PIN_XY=14322,-7874,14292,-7933,14262,-7874 $DEVICE_ID=1001
MM425 34 54 119 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13956 $Y=-6809  $PIN_XY=13986,-6726,13956,-6809,13926,-6726 $DEVICE_ID=1001
MM426 34 53 87 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13956 $Y=-7933  $PIN_XY=13986,-7874,13956,-7933,13926,-7874 $DEVICE_ID=1001
MM427 GND! 120 119 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13620 $Y=-6457  $PIN_XY=(13650,-6552,13650,-6726),13620,-6457,(13590,-6552,13590,-6726) $DEVICE_ID=1001
MM428 GND! 88 87 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13620 $Y=-7596  $PIN_XY=(13650,-7700,13650,-7874),13620,-7596,(13590,-7700,13590,-7874) $DEVICE_ID=1001
MM429 120 119 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13284 $Y=-6457  $PIN_XY=(13314,-6552,13314,-6726),13284,-6457,(13254,-6552,13254,-6726) $DEVICE_ID=1001
MM430 88 87 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=13284 $Y=-7581  $PIN_XY=(13314,-7700,13314,-7874),13284,-7581,(13254,-7700,13254,-7874) $DEVICE_ID=1001
MM431 120 54 33 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12948 $Y=-6809  $PIN_XY=12978,-6726,12948,-6809,12918,-6726 $DEVICE_ID=1001
MM432 88 53 33 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12948 $Y=-7933  $PIN_XY=12978,-7874,12948,-7933,12918,-7874 $DEVICE_ID=1001
MM433 32 54 117 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12612 $Y=-6809  $PIN_XY=12642,-6726,12612,-6809,12582,-6726 $DEVICE_ID=1001
MM434 32 53 85 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12612 $Y=-7933  $PIN_XY=12642,-7874,12612,-7933,12582,-7874 $DEVICE_ID=1001
MM435 GND! 118 117 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=12276 $Y=-6457  $PIN_XY=(12306,-6552,12306,-6726),12276,-6457,(12246,-6552,12246,-6726) $DEVICE_ID=1001
MM436 GND! 86 85 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=12276 $Y=-7581  $PIN_XY=(12306,-7700,12306,-7874),12276,-7581,(12246,-7700,12246,-7874) $DEVICE_ID=1001
MM437 118 117 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11940 $Y=-6457  $PIN_XY=(11970,-6552,11970,-6726),11940,-6457,(11910,-6552,11910,-6726) $DEVICE_ID=1001
MM438 86 85 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=11940 $Y=-7581  $PIN_XY=(11970,-7700,11970,-7874),11940,-7581,(11910,-7700,11910,-7874) $DEVICE_ID=1001
MM439 118 54 31 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11604 $Y=-6809  $PIN_XY=11634,-6726,11604,-6809,11574,-6726 $DEVICE_ID=1001
MM440 86 53 31 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11604 $Y=-7933  $PIN_XY=11634,-7874,11604,-7933,11574,-7874 $DEVICE_ID=1001
MM441 30 54 115 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11268 $Y=-6809  $PIN_XY=11298,-6726,11268,-6809,11238,-6726 $DEVICE_ID=1001
MM442 30 53 83 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11268 $Y=-7933  $PIN_XY=11298,-7874,11268,-7933,11238,-7874 $DEVICE_ID=1001
MM443 GND! 116 115 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10932 $Y=-6457  $PIN_XY=(10962,-6552,10962,-6726),10932,-6457,(10902,-6552,10902,-6726) $DEVICE_ID=1001
MM444 GND! 84 83 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10932 $Y=-7581  $PIN_XY=(10962,-7700,10962,-7874),10932,-7581,(10902,-7700,10902,-7874) $DEVICE_ID=1001
MM445 116 115 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10596 $Y=-6457  $PIN_XY=(10626,-6552,10626,-6726),10596,-6457,(10566,-6552,10566,-6726) $DEVICE_ID=1001
MM446 84 83 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=10596 $Y=-7581  $PIN_XY=(10626,-7700,10626,-7874),10596,-7581,(10566,-7700,10566,-7874) $DEVICE_ID=1001
MM447 116 54 29 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10260 $Y=-6809  $PIN_XY=10290,-6726,10260,-6809,10230,-6726 $DEVICE_ID=1001
MM448 84 53 29 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10260 $Y=-7933  $PIN_XY=10290,-7874,10260,-7933,10230,-7874 $DEVICE_ID=1001
MM449 28 54 113 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9924 $Y=-6809  $PIN_XY=9954,-6726,9924,-6809,9894,-6726 $DEVICE_ID=1001
MM450 28 53 81 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9924 $Y=-7933  $PIN_XY=9954,-7874,9924,-7933,9894,-7874 $DEVICE_ID=1001
MM451 GND! 114 113 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9588 $Y=-6457  $PIN_XY=(9618,-6552,9618,-6726),9588,-6457,(9558,-6552,9558,-6726) $DEVICE_ID=1001
MM452 GND! 82 81 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9588 $Y=-7581  $PIN_XY=(9618,-7700,9618,-7874),9588,-7581,(9558,-7700,9558,-7874) $DEVICE_ID=1001
MM453 114 113 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9252 $Y=-6457  $PIN_XY=(9282,-6552,9282,-6726),9252,-6457,(9222,-6552,9222,-6726) $DEVICE_ID=1001
MM454 82 81 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=9252 $Y=-7581  $PIN_XY=(9282,-7700,9282,-7874),9252,-7581,(9222,-7700,9222,-7874) $DEVICE_ID=1001
MM455 114 54 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8916 $Y=-6809  $PIN_XY=8946,-6726,8916,-6809,8886,-6726 $DEVICE_ID=1001
MM456 82 53 27 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8916 $Y=-7933  $PIN_XY=8946,-7874,8916,-7933,8886,-7874 $DEVICE_ID=1001
MM457 26 54 111 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8580 $Y=-6809  $PIN_XY=8610,-6726,8580,-6809,8550,-6726 $DEVICE_ID=1001
MM458 26 53 79 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8580 $Y=-7933  $PIN_XY=8610,-7874,8580,-7933,8550,-7874 $DEVICE_ID=1001
MM459 GND! 112 111 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8244 $Y=-6457  $PIN_XY=(8274,-6552,8274,-6726),8244,-6457,(8214,-6552,8214,-6726) $DEVICE_ID=1001
MM460 GND! 80 79 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=8244 $Y=-7581  $PIN_XY=(8274,-7700,8274,-7874),8244,-7581,(8214,-7700,8214,-7874) $DEVICE_ID=1001
MM461 112 111 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7908 $Y=-6457  $PIN_XY=(7938,-6552,7938,-6726),7908,-6457,(7878,-6552,7878,-6726) $DEVICE_ID=1001
MM462 80 79 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=7908 $Y=-7581  $PIN_XY=(7938,-7700,7938,-7874),7908,-7581,(7878,-7700,7878,-7874) $DEVICE_ID=1001
MM463 112 54 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7572 $Y=-6809  $PIN_XY=7602,-6726,7572,-6809,7542,-6726 $DEVICE_ID=1001
MM464 80 53 25 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7572 $Y=-7933  $PIN_XY=7602,-7874,7572,-7933,7542,-7874 $DEVICE_ID=1001
MM465 24 54 109 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7236 $Y=-6809  $PIN_XY=7266,-6726,7236,-6809,7206,-6726 $DEVICE_ID=1001
MM466 24 53 77 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7236 $Y=-7933  $PIN_XY=7266,-7874,7236,-7933,7206,-7874 $DEVICE_ID=1001
MM467 GND! 110 109 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6900 $Y=-6457  $PIN_XY=(6930,-6552,6930,-6726),6900,-6457,(6870,-6552,6870,-6726) $DEVICE_ID=1001
MM468 GND! 78 77 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6900 $Y=-7581  $PIN_XY=(6930,-7700,6930,-7874),6900,-7581,(6870,-7700,6870,-7874) $DEVICE_ID=1001
MM469 110 109 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6564 $Y=-6457  $PIN_XY=(6594,-6552,6594,-6726),6564,-6457,(6534,-6552,6534,-6726) $DEVICE_ID=1001
MM470 78 77 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=6564 $Y=-7581  $PIN_XY=(6594,-7700,6594,-7874),6564,-7581,(6534,-7700,6534,-7874) $DEVICE_ID=1001
MM471 110 54 23 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6228 $Y=-6809  $PIN_XY=6258,-6726,6228,-6809,6198,-6726 $DEVICE_ID=1001
MM472 78 53 23 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6228 $Y=-7933  $PIN_XY=6258,-7874,6228,-7933,6198,-7874 $DEVICE_ID=1001
MM473 22 54 107 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5892 $Y=-6809  $PIN_XY=5922,-6726,5892,-6809,5862,-6726 $DEVICE_ID=1001
MM474 22 53 75 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5892 $Y=-7933  $PIN_XY=5922,-7874,5892,-7933,5862,-7874 $DEVICE_ID=1001
MM475 GND! 108 107 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5556 $Y=-6457  $PIN_XY=(5586,-6552,5586,-6726),5556,-6457,(5526,-6552,5526,-6726) $DEVICE_ID=1001
MM476 GND! 76 75 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5556 $Y=-7581  $PIN_XY=(5586,-7700,5586,-7874),5556,-7581,(5526,-7700,5526,-7874) $DEVICE_ID=1001
MM477 108 107 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5220 $Y=-6457  $PIN_XY=(5250,-6552,5250,-6726),5220,-6457,(5190,-6552,5190,-6726) $DEVICE_ID=1001
MM478 76 75 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=5220 $Y=-7581  $PIN_XY=(5250,-7700,5250,-7874),5220,-7581,(5190,-7700,5190,-7874) $DEVICE_ID=1001
MM479 108 54 21 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4884 $Y=-6809  $PIN_XY=4914,-6726,4884,-6809,4854,-6726 $DEVICE_ID=1001
MM480 76 53 21 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4884 $Y=-7933  $PIN_XY=4914,-7874,4884,-7933,4854,-7874 $DEVICE_ID=1001
MM481 20 54 105 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4548 $Y=-6809  $PIN_XY=4578,-6726,4548,-6809,4518,-6726 $DEVICE_ID=1001
MM482 20 53 73 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4548 $Y=-7933  $PIN_XY=4578,-7874,4548,-7933,4518,-7874 $DEVICE_ID=1001
MM483 GND! 106 105 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4212 $Y=-6457  $PIN_XY=(4242,-6552,4242,-6726),4212,-6457,(4182,-6552,4182,-6726) $DEVICE_ID=1001
MM484 GND! 74 73 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=4212 $Y=-7581  $PIN_XY=(4242,-7700,4242,-7874),4212,-7581,(4182,-7700,4182,-7874) $DEVICE_ID=1001
MM485 106 105 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3876 $Y=-6457  $PIN_XY=(3906,-6552,3906,-6726),3876,-6457,(3846,-6552,3846,-6726) $DEVICE_ID=1001
MM486 74 73 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=3876 $Y=-7581  $PIN_XY=(3906,-7700,3906,-7874),3876,-7581,(3846,-7700,3846,-7874) $DEVICE_ID=1001
MM487 106 54 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3540 $Y=-6809  $PIN_XY=3570,-6726,3540,-6809,3510,-6726 $DEVICE_ID=1001
MM488 74 53 19 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3540 $Y=-7933  $PIN_XY=3570,-7874,3540,-7933,3510,-7874 $DEVICE_ID=1001
MM489 18 54 103 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3204 $Y=-6809  $PIN_XY=3234,-6726,3204,-6809,3174,-6726 $DEVICE_ID=1001
MM490 18 53 71 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3204 $Y=-7933  $PIN_XY=3234,-7874,3204,-7933,3174,-7874 $DEVICE_ID=1001
MM491 GND! 104 103 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2868 $Y=-6457  $PIN_XY=(2898,-6552,2898,-6726),2868,-6457,(2838,-6552,2838,-6726) $DEVICE_ID=1001
MM492 GND! 72 71 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2868 $Y=-7581  $PIN_XY=(2898,-7700,2898,-7874),2868,-7581,(2838,-7700,2838,-7874) $DEVICE_ID=1001
MM493 104 103 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2532 $Y=-6457  $PIN_XY=(2562,-6552,2562,-6726),2532,-6457,(2502,-6552,2502,-6726) $DEVICE_ID=1001
MM494 72 71 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=2532 $Y=-7581  $PIN_XY=(2562,-7700,2562,-7874),2532,-7581,(2502,-7700,2502,-7874) $DEVICE_ID=1001
MM495 104 54 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2196 $Y=-6809  $PIN_XY=2226,-6726,2196,-6809,2166,-6726 $DEVICE_ID=1001
MM496 72 53 17 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2196 $Y=-7933  $PIN_XY=2226,-7874,2196,-7933,2166,-7874 $DEVICE_ID=1001
MM497 16 54 101 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1860 $Y=-6809  $PIN_XY=1890,-6726,1860,-6809,1830,-6726 $DEVICE_ID=1001
MM498 16 53 69 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1860 $Y=-7933  $PIN_XY=1890,-7874,1860,-7933,1830,-7874 $DEVICE_ID=1001
MM499 GND! 102 101 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1524 $Y=-6457  $PIN_XY=(1554,-6552,1554,-6726),1524,-6457,(1494,-6552,1494,-6726) $DEVICE_ID=1001
MM500 GND! 70 69 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1524 $Y=-7581  $PIN_XY=(1554,-7700,1554,-7874),1524,-7581,(1494,-7700,1494,-7874) $DEVICE_ID=1001
MM501 102 101 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1188 $Y=-6457  $PIN_XY=(1218,-6552,1218,-6726),1188,-6457,(1158,-6552,1158,-6726) $DEVICE_ID=1001
MM502 70 69 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=1188 $Y=-7581  $PIN_XY=(1218,-7700,1218,-7874),1188,-7581,(1158,-7700,1158,-7874) $DEVICE_ID=1001
MM503 102 54 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=852 $Y=-6809  $PIN_XY=882,-6726,852,-6809,822,-6726 $DEVICE_ID=1001
MM504 70 53 15 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=852 $Y=-7933  $PIN_XY=882,-7874,852,-7933,822,-7874 $DEVICE_ID=1001
MM505 13 54 99 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=516 $Y=-6809  $PIN_XY=546,-6726,516,-6809,486,-6726 $DEVICE_ID=1001
MM506 13 53 67 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=516 $Y=-7933  $PIN_XY=546,-7874,516,-7933,486,-7874 $DEVICE_ID=1001
MM507 GND! 100 99 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=180 $Y=-6457  $PIN_XY=(210,-6552,210,-6726),180,-6457,(150,-6552,150,-6726) $DEVICE_ID=1001
MM508 GND! 68 67 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=180 $Y=-7581  $PIN_XY=(210,-7700,210,-7874),180,-7581,(150,-7700,150,-7874) $DEVICE_ID=1001
MM509 100 99 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=-156 $Y=-6457  $PIN_XY=(-126,-6552,-126,-6726),-156,-6457,(-186,-6552,-186,-6726) $DEVICE_ID=1001
MM510 68 67 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=-156 $Y=-7581  $PIN_XY=(-126,-7700,-126,-7874),-156,-7581,(-186,-7700,-186,-7874) $DEVICE_ID=1001
MM511 100 54 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=-492 $Y=-6809  $PIN_XY=-462,-6726,-492,-6809,-522,-6726 $DEVICE_ID=1001
MM512 68 53 12 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=-492 $Y=-7933  $PIN_XY=-462,-7874,-492,-7933,-522,-7874 $DEVICE_ID=1001
MM513 Q<0> 334 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=24374 $Y=-20862  $PIN_XY=24404,-21038,24374,-20862,24344,-21038 $DEVICE_ID=1001
MM514 Q<1> 330 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=24374 $Y=-22750  $PIN_XY=24404,-22926,24374,-22750,24344,-22926 $DEVICE_ID=1001
MM515 334 333 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=24038 $Y=-20863  $PIN_XY=24068,-21038,24038,-20863,24008,-21038 $DEVICE_ID=1001
MM516 330 329 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=24038 $Y=-22751  $PIN_XY=24068,-22926,24038,-22751,24008,-22926 $DEVICE_ID=1001
MM517 333 CLK 1544 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=23702 $Y=-21209  $PIN_XY=23732,-21208,23702,-21209,23672,-21208 $DEVICE_ID=1001
MM518 329 CLK 1542 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=23702 $Y=-23097  $PIN_XY=23732,-23096,23702,-23097,23672,-23096 $DEVICE_ID=1001
MM519 1544 332 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=23534 $Y=-21216  $PIN_XY=23564,-21208,23534,-21216,23504,-21208 $DEVICE_ID=1001
MM520 1542 328 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=23534 $Y=-23104  $PIN_XY=23564,-23096,23534,-23104,23504,-23096 $DEVICE_ID=1001
MM521 332 331 1543 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=23198 $Y=-21141  $PIN_XY=(23228,-21038,23228,-21208),23198,-21141,(23168,-21038,23168,-21208) $DEVICE_ID=1001
MM522 328 327 1541 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=23198 $Y=-23029  $PIN_XY=(23228,-22926,23228,-23096),23198,-23029,(23168,-22926,23168,-23096) $DEVICE_ID=1001
MM523 1543 CLK GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=23030 $Y=-21124  $PIN_XY=(23060,-21038,23060,-21208),23030,-21124,(23000,-21038,23000,-21208) $DEVICE_ID=1001
MM524 1541 CLK GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=23030 $Y=-23012  $PIN_XY=(23060,-22926,23060,-23096),23030,-23012,(23000,-22926,23000,-23096) $DEVICE_ID=1001
MM525 331 2 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=22694 $Y=-21210  $PIN_XY=22724,-21208,22694,-21210,22664,-21208 $DEVICE_ID=1001
MM526 327 4 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=22694 $Y=-23098  $PIN_XY=22724,-23096,22694,-23098,22664,-23096 $DEVICE_ID=1001
MM527 Q<2> 338 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=24374 $Y=-24638  $PIN_XY=24404,-24814,24374,-24638,24344,-24814 $DEVICE_ID=1001
MM528 Q<3> 326 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=24374 $Y=-26526  $PIN_XY=24404,-26702,24374,-26526,24344,-26702 $DEVICE_ID=1001
MM529 338 337 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=24038 $Y=-24639  $PIN_XY=24068,-24814,24038,-24639,24008,-24814 $DEVICE_ID=1001
MM530 326 325 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=24038 $Y=-26527  $PIN_XY=24068,-26702,24038,-26527,24008,-26702 $DEVICE_ID=1001
MM531 337 CLK 1546 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=23702 $Y=-24985  $PIN_XY=23732,-24984,23702,-24985,23672,-24984 $DEVICE_ID=1001
MM532 325 CLK 1540 nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=23702 $Y=-26873  $PIN_XY=23732,-26872,23702,-26873,23672,-26872 $DEVICE_ID=1001
MM533 1546 336 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=23534 $Y=-24992  $PIN_XY=23564,-24984,23534,-24992,23504,-24984 $DEVICE_ID=1001
MM534 1540 324 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=23534 $Y=-26880  $PIN_XY=23564,-26872,23534,-26880,23504,-26872 $DEVICE_ID=1001
MM535 336 335 1545 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=23198 $Y=-24917  $PIN_XY=(23228,-24814,23228,-24984),23198,-24917,(23168,-24814,23168,-24984) $DEVICE_ID=1001
MM536 324 323 1539 nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=1.134e-15 PDEO=1.17e-07
+	 PSEO=2.34e-07 $X=23198 $Y=-26805  $PIN_XY=(23228,-26702,23228,-26872),23198,-26805,(23168,-26702,23168,-26872) $DEVICE_ID=1001
MM537 1545 CLK GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=23030 $Y=-24900  $PIN_XY=(23060,-24814,23060,-24984),23030,-24900,(23000,-24814,23000,-24984) $DEVICE_ID=1001
MM538 1539 CLK GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=1.134e-15 ASEO=5.67e-16 PDEO=2.34e-07
+	 PSEO=1.17e-07 $X=23030 $Y=-26788  $PIN_XY=(23060,-26702,23060,-26872),23030,-26788,(23000,-26702,23000,-26872) $DEVICE_ID=1001
MM539 335 8 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=22694 $Y=-24986  $PIN_XY=22724,-24984,22694,-24986,22664,-24984 $DEVICE_ID=1001
MM540 323 6 GND! nmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=22694 $Y=-26874  $PIN_XY=22724,-26872,22694,-26874,22664,-26872 $DEVICE_ID=1001
MM541 VDD! 322 321 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20340 $Y=304  $PIN_XY=20370,502,20340,304,20310,502 $DEVICE_ID=1003
MM542 VDD! 290 289 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20340 $Y=-720  $PIN_XY=20370,-646,20340,-720,20310,-646 $DEVICE_ID=1003
MM543 VDD! 258 257 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20340 $Y=-1867  $PIN_XY=20370,-1792,20340,-1867,20310,-1792 $DEVICE_ID=1003
MM544 322 321 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20004 $Y=304  $PIN_XY=20034,502,20004,304,19974,502 $DEVICE_ID=1003
MM545 290 289 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20004 $Y=-720  $PIN_XY=20034,-646,20004,-720,19974,-646 $DEVICE_ID=1003
MM546 258 257 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20004 $Y=-1867  $PIN_XY=20034,-1792,20004,-1867,19974,-1792 $DEVICE_ID=1003
MM547 VDD! 320 319 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18996 $Y=304  $PIN_XY=19026,502,18996,304,18966,502 $DEVICE_ID=1003
MM548 VDD! 288 287 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18996 $Y=-720  $PIN_XY=19026,-646,18996,-720,18966,-646 $DEVICE_ID=1003
MM549 VDD! 256 255 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18996 $Y=-1867  $PIN_XY=19026,-1792,18996,-1867,18966,-1792 $DEVICE_ID=1003
MM550 320 319 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18660 $Y=304  $PIN_XY=18690,502,18660,304,18630,502 $DEVICE_ID=1003
MM551 288 287 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18660 $Y=-720  $PIN_XY=18690,-646,18660,-720,18630,-646 $DEVICE_ID=1003
MM552 256 255 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18660 $Y=-1867  $PIN_XY=18690,-1792,18660,-1867,18630,-1792 $DEVICE_ID=1003
MM553 VDD! 318 317 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17652 $Y=304  $PIN_XY=17682,502,17652,304,17622,502 $DEVICE_ID=1003
MM554 VDD! 286 285 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17652 $Y=-720  $PIN_XY=17682,-646,17652,-720,17622,-646 $DEVICE_ID=1003
MM555 VDD! 254 253 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17652 $Y=-1867  $PIN_XY=17682,-1792,17652,-1867,17622,-1792 $DEVICE_ID=1003
MM556 318 317 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17316 $Y=304  $PIN_XY=17346,502,17316,304,17286,502 $DEVICE_ID=1003
MM557 286 285 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17316 $Y=-720  $PIN_XY=17346,-646,17316,-720,17286,-646 $DEVICE_ID=1003
MM558 254 253 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17316 $Y=-1867  $PIN_XY=17346,-1792,17316,-1867,17286,-1792 $DEVICE_ID=1003
MM559 VDD! 316 315 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16308 $Y=304  $PIN_XY=16338,502,16308,304,16278,502 $DEVICE_ID=1003
MM560 VDD! 284 283 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16308 $Y=-720  $PIN_XY=16338,-646,16308,-720,16278,-646 $DEVICE_ID=1003
MM561 VDD! 252 251 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16308 $Y=-1867  $PIN_XY=16338,-1792,16308,-1867,16278,-1792 $DEVICE_ID=1003
MM562 316 315 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15972 $Y=304  $PIN_XY=16002,502,15972,304,15942,502 $DEVICE_ID=1003
MM563 284 283 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15972 $Y=-720  $PIN_XY=16002,-646,15972,-720,15942,-646 $DEVICE_ID=1003
MM564 252 251 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15972 $Y=-1867  $PIN_XY=16002,-1792,15972,-1867,15942,-1792 $DEVICE_ID=1003
MM565 VDD! 314 313 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14964 $Y=304  $PIN_XY=14994,502,14964,304,14934,502 $DEVICE_ID=1003
MM566 VDD! 282 281 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14964 $Y=-720  $PIN_XY=14994,-646,14964,-720,14934,-646 $DEVICE_ID=1003
MM567 VDD! 250 249 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14964 $Y=-1867  $PIN_XY=14994,-1792,14964,-1867,14934,-1792 $DEVICE_ID=1003
MM568 314 313 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14628 $Y=304  $PIN_XY=14658,502,14628,304,14598,502 $DEVICE_ID=1003
MM569 282 281 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14628 $Y=-720  $PIN_XY=14658,-646,14628,-720,14598,-646 $DEVICE_ID=1003
MM570 VDD! 312 311 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13620 $Y=304  $PIN_XY=13650,502,13620,304,13590,502 $DEVICE_ID=1003
MM571 VDD! 280 279 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13620 $Y=-720  $PIN_XY=13650,-646,13620,-720,13590,-646 $DEVICE_ID=1003
MM572 312 311 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13284 $Y=304  $PIN_XY=13314,502,13284,304,13254,502 $DEVICE_ID=1003
MM573 280 279 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13284 $Y=-720  $PIN_XY=13314,-646,13284,-720,13254,-646 $DEVICE_ID=1003
MM574 250 249 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14628 $Y=-1867  $PIN_XY=14658,-1792,14628,-1867,14598,-1792 $DEVICE_ID=1003
MM575 VDD! 248 247 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13620 $Y=-1867  $PIN_XY=13650,-1792,13620,-1867,13590,-1792 $DEVICE_ID=1003
MM576 248 247 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13284 $Y=-1867  $PIN_XY=13314,-1792,13284,-1867,13254,-1792 $DEVICE_ID=1003
MM577 VDD! 310 309 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12276 $Y=304  $PIN_XY=12306,502,12276,304,12246,502 $DEVICE_ID=1003
MM578 VDD! 278 277 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12276 $Y=-720  $PIN_XY=12306,-646,12276,-720,12246,-646 $DEVICE_ID=1003
MM579 VDD! 246 245 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12276 $Y=-1867  $PIN_XY=12306,-1792,12276,-1867,12246,-1792 $DEVICE_ID=1003
MM580 310 309 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11940 $Y=304  $PIN_XY=11970,502,11940,304,11910,502 $DEVICE_ID=1003
MM581 278 277 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11940 $Y=-720  $PIN_XY=11970,-646,11940,-720,11910,-646 $DEVICE_ID=1003
MM582 246 245 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11940 $Y=-1867  $PIN_XY=11970,-1792,11940,-1867,11910,-1792 $DEVICE_ID=1003
MM583 VDD! 308 307 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10932 $Y=304  $PIN_XY=10962,502,10932,304,10902,502 $DEVICE_ID=1003
MM584 VDD! 276 275 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10932 $Y=-720  $PIN_XY=10962,-646,10932,-720,10902,-646 $DEVICE_ID=1003
MM585 VDD! 244 243 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10932 $Y=-1867  $PIN_XY=10962,-1792,10932,-1867,10902,-1792 $DEVICE_ID=1003
MM586 308 307 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10596 $Y=304  $PIN_XY=10626,502,10596,304,10566,502 $DEVICE_ID=1003
MM587 VDD! 306 305 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9588 $Y=304  $PIN_XY=9618,502,9588,304,9558,502 $DEVICE_ID=1003
MM588 306 305 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9252 $Y=304  $PIN_XY=9282,502,9252,304,9222,502 $DEVICE_ID=1003
MM589 276 275 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10596 $Y=-720  $PIN_XY=10626,-646,10596,-720,10566,-646 $DEVICE_ID=1003
MM590 244 243 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10596 $Y=-1867  $PIN_XY=10626,-1792,10596,-1867,10566,-1792 $DEVICE_ID=1003
MM591 VDD! 274 273 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9588 $Y=-720  $PIN_XY=9618,-646,9588,-720,9558,-646 $DEVICE_ID=1003
MM592 VDD! 242 241 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9588 $Y=-1867  $PIN_XY=9618,-1792,9588,-1867,9558,-1792 $DEVICE_ID=1003
MM593 274 273 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9252 $Y=-720  $PIN_XY=9282,-646,9252,-720,9222,-646 $DEVICE_ID=1003
MM594 242 241 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9252 $Y=-1867  $PIN_XY=9282,-1792,9252,-1867,9222,-1792 $DEVICE_ID=1003
MM595 VDD! 304 303 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8244 $Y=304  $PIN_XY=8274,502,8244,304,8214,502 $DEVICE_ID=1003
MM596 VDD! 272 271 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8244 $Y=-720  $PIN_XY=8274,-646,8244,-720,8214,-646 $DEVICE_ID=1003
MM597 304 303 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7908 $Y=304  $PIN_XY=7938,502,7908,304,7878,502 $DEVICE_ID=1003
MM598 272 271 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7908 $Y=-720  $PIN_XY=7938,-646,7908,-720,7878,-646 $DEVICE_ID=1003
MM599 VDD! 302 301 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6900 $Y=304  $PIN_XY=6930,502,6900,304,6870,502 $DEVICE_ID=1003
MM600 VDD! 270 269 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6900 $Y=-720  $PIN_XY=6930,-646,6900,-720,6870,-646 $DEVICE_ID=1003
MM601 VDD! 240 239 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8244 $Y=-1867  $PIN_XY=8274,-1792,8244,-1867,8214,-1792 $DEVICE_ID=1003
MM602 240 239 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7908 $Y=-1867  $PIN_XY=7938,-1792,7908,-1867,7878,-1792 $DEVICE_ID=1003
MM603 VDD! 238 237 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6900 $Y=-1867  $PIN_XY=6930,-1792,6900,-1867,6870,-1792 $DEVICE_ID=1003
MM604 302 301 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6564 $Y=304  $PIN_XY=6594,502,6564,304,6534,502 $DEVICE_ID=1003
MM605 270 269 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6564 $Y=-720  $PIN_XY=6594,-646,6564,-720,6534,-646 $DEVICE_ID=1003
MM606 238 237 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6564 $Y=-1867  $PIN_XY=6594,-1792,6564,-1867,6534,-1792 $DEVICE_ID=1003
MM607 VDD! 300 299 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5556 $Y=304  $PIN_XY=5586,502,5556,304,5526,502 $DEVICE_ID=1003
MM608 VDD! 268 267 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5556 $Y=-720  $PIN_XY=5586,-646,5556,-720,5526,-646 $DEVICE_ID=1003
MM609 VDD! 236 235 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5556 $Y=-1867  $PIN_XY=5586,-1792,5556,-1867,5526,-1792 $DEVICE_ID=1003
MM610 300 299 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5220 $Y=304  $PIN_XY=5250,502,5220,304,5190,502 $DEVICE_ID=1003
MM611 268 267 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5220 $Y=-720  $PIN_XY=5250,-646,5220,-720,5190,-646 $DEVICE_ID=1003
MM612 236 235 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5220 $Y=-1867  $PIN_XY=5250,-1792,5220,-1867,5190,-1792 $DEVICE_ID=1003
MM613 VDD! 298 297 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4212 $Y=304  $PIN_XY=4242,502,4212,304,4182,502 $DEVICE_ID=1003
MM614 VDD! 266 265 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4212 $Y=-720  $PIN_XY=4242,-646,4212,-720,4182,-646 $DEVICE_ID=1003
MM615 VDD! 234 233 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4212 $Y=-1867  $PIN_XY=4242,-1792,4212,-1867,4182,-1792 $DEVICE_ID=1003
MM616 298 297 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3876 $Y=304  $PIN_XY=3906,502,3876,304,3846,502 $DEVICE_ID=1003
MM617 266 265 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3876 $Y=-720  $PIN_XY=3906,-646,3876,-720,3846,-646 $DEVICE_ID=1003
MM618 234 233 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3876 $Y=-1867  $PIN_XY=3906,-1792,3876,-1867,3846,-1792 $DEVICE_ID=1003
MM619 VDD! 296 295 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2868 $Y=304  $PIN_XY=2898,502,2868,304,2838,502 $DEVICE_ID=1003
MM620 VDD! 264 263 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2868 $Y=-720  $PIN_XY=2898,-646,2868,-720,2838,-646 $DEVICE_ID=1003
MM621 VDD! 232 231 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2868 $Y=-1867  $PIN_XY=2898,-1792,2868,-1867,2838,-1792 $DEVICE_ID=1003
MM622 296 295 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2532 $Y=304  $PIN_XY=2562,502,2532,304,2502,502 $DEVICE_ID=1003
MM623 264 263 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2532 $Y=-720  $PIN_XY=2562,-646,2532,-720,2502,-646 $DEVICE_ID=1003
MM624 232 231 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2532 $Y=-1867  $PIN_XY=2562,-1792,2532,-1867,2502,-1792 $DEVICE_ID=1003
MM625 VDD! 294 293 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1524 $Y=304  $PIN_XY=1554,502,1524,304,1494,502 $DEVICE_ID=1003
MM626 VDD! 262 261 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1524 $Y=-720  $PIN_XY=1554,-646,1524,-720,1494,-646 $DEVICE_ID=1003
MM627 VDD! 230 229 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1524 $Y=-1867  $PIN_XY=1554,-1792,1524,-1867,1494,-1792 $DEVICE_ID=1003
MM628 294 293 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1188 $Y=304  $PIN_XY=1218,502,1188,304,1158,502 $DEVICE_ID=1003
MM629 262 261 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1188 $Y=-720  $PIN_XY=1218,-646,1188,-720,1158,-646 $DEVICE_ID=1003
MM630 230 229 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1188 $Y=-1867  $PIN_XY=1218,-1792,1188,-1867,1158,-1792 $DEVICE_ID=1003
MM631 VDD! 292 291 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=180 $Y=304  $PIN_XY=210,502,180,304,150,502 $DEVICE_ID=1003
MM632 VDD! 260 259 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=180 $Y=-720  $PIN_XY=210,-646,180,-720,150,-646 $DEVICE_ID=1003
MM633 VDD! 228 227 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=180 $Y=-1867  $PIN_XY=210,-1792,180,-1867,150,-1792 $DEVICE_ID=1003
MM634 292 291 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=-156 $Y=304  $PIN_XY=-126,502,-156,304,-186,502 $DEVICE_ID=1003
MM635 260 259 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=-156 $Y=-720  $PIN_XY=-126,-646,-156,-720,-186,-646 $DEVICE_ID=1003
MM636 228 227 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=-156 $Y=-1867  $PIN_XY=-126,-1792,-156,-1867,-186,-1792 $DEVICE_ID=1003
MM637 VDD! 226 225 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20340 $Y=-3012  $PIN_XY=20370,-2940,20340,-3012,20310,-2940 $DEVICE_ID=1003
MM638 VDD! 194 193 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20340 $Y=-4160  $PIN_XY=20370,-4088,20340,-4160,20310,-4088 $DEVICE_ID=1003
MM639 VDD! 162 161 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20340 $Y=-5310  $PIN_XY=20370,-5236,20340,-5310,20310,-5236 $DEVICE_ID=1003
MM640 226 225 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20004 $Y=-3012  $PIN_XY=20034,-2940,20004,-3012,19974,-2940 $DEVICE_ID=1003
MM641 194 193 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20004 $Y=-4160  $PIN_XY=20034,-4088,20004,-4160,19974,-4088 $DEVICE_ID=1003
MM642 162 161 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20004 $Y=-5310  $PIN_XY=20034,-5236,20004,-5310,19974,-5236 $DEVICE_ID=1003
MM643 VDD! 224 223 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18996 $Y=-3012  $PIN_XY=19026,-2940,18996,-3012,18966,-2940 $DEVICE_ID=1003
MM644 VDD! 192 191 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18996 $Y=-4160  $PIN_XY=19026,-4088,18996,-4160,18966,-4088 $DEVICE_ID=1003
MM645 VDD! 160 159 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18996 $Y=-5310  $PIN_XY=19026,-5236,18996,-5310,18966,-5236 $DEVICE_ID=1003
MM646 224 223 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18660 $Y=-3012  $PIN_XY=18690,-2940,18660,-3012,18630,-2940 $DEVICE_ID=1003
MM647 192 191 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18660 $Y=-4160  $PIN_XY=18690,-4088,18660,-4160,18630,-4088 $DEVICE_ID=1003
MM648 160 159 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18660 $Y=-5310  $PIN_XY=18690,-5236,18660,-5310,18630,-5236 $DEVICE_ID=1003
MM649 VDD! 222 221 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17652 $Y=-3012  $PIN_XY=17682,-2940,17652,-3012,17622,-2940 $DEVICE_ID=1003
MM650 VDD! 190 189 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17652 $Y=-4160  $PIN_XY=17682,-4088,17652,-4160,17622,-4088 $DEVICE_ID=1003
MM651 VDD! 158 157 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17652 $Y=-5310  $PIN_XY=17682,-5236,17652,-5310,17622,-5236 $DEVICE_ID=1003
MM652 222 221 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17316 $Y=-3012  $PIN_XY=17346,-2940,17316,-3012,17286,-2940 $DEVICE_ID=1003
MM653 190 189 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17316 $Y=-4160  $PIN_XY=17346,-4088,17316,-4160,17286,-4088 $DEVICE_ID=1003
MM654 158 157 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17316 $Y=-5310  $PIN_XY=17346,-5236,17316,-5310,17286,-5236 $DEVICE_ID=1003
MM655 VDD! 220 219 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16308 $Y=-3012  $PIN_XY=16338,-2940,16308,-3012,16278,-2940 $DEVICE_ID=1003
MM656 VDD! 188 187 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16308 $Y=-4160  $PIN_XY=16338,-4088,16308,-4160,16278,-4088 $DEVICE_ID=1003
MM657 VDD! 156 155 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16308 $Y=-5310  $PIN_XY=16338,-5236,16308,-5310,16278,-5236 $DEVICE_ID=1003
MM658 220 219 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15972 $Y=-3012  $PIN_XY=16002,-2940,15972,-3012,15942,-2940 $DEVICE_ID=1003
MM659 188 187 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15972 $Y=-4160  $PIN_XY=16002,-4088,15972,-4160,15942,-4088 $DEVICE_ID=1003
MM660 156 155 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15972 $Y=-5310  $PIN_XY=16002,-5236,15972,-5310,15942,-5236 $DEVICE_ID=1003
MM661 VDD! 218 217 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14964 $Y=-3012  $PIN_XY=14994,-2940,14964,-3012,14934,-2940 $DEVICE_ID=1003
MM662 VDD! 186 185 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14964 $Y=-4160  $PIN_XY=14994,-4088,14964,-4160,14934,-4088 $DEVICE_ID=1003
MM663 VDD! 154 153 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14964 $Y=-5310  $PIN_XY=14994,-5236,14964,-5310,14934,-5236 $DEVICE_ID=1003
MM664 218 217 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14628 $Y=-3012  $PIN_XY=14658,-2940,14628,-3012,14598,-2940 $DEVICE_ID=1003
MM665 186 185 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14628 $Y=-4160  $PIN_XY=14658,-4088,14628,-4160,14598,-4088 $DEVICE_ID=1003
MM666 154 153 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14628 $Y=-5310  $PIN_XY=14658,-5236,14628,-5310,14598,-5236 $DEVICE_ID=1003
MM667 VDD! 216 215 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13620 $Y=-3012  $PIN_XY=13650,-2940,13620,-3012,13590,-2940 $DEVICE_ID=1003
MM668 VDD! 184 183 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13620 $Y=-4160  $PIN_XY=13650,-4088,13620,-4160,13590,-4088 $DEVICE_ID=1003
MM669 VDD! 152 151 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13620 $Y=-5310  $PIN_XY=13650,-5236,13620,-5310,13590,-5236 $DEVICE_ID=1003
MM670 216 215 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13284 $Y=-3012  $PIN_XY=13314,-2940,13284,-3012,13254,-2940 $DEVICE_ID=1003
MM671 184 183 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13284 $Y=-4160  $PIN_XY=13314,-4088,13284,-4160,13254,-4088 $DEVICE_ID=1003
MM672 152 151 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13284 $Y=-5310  $PIN_XY=13314,-5236,13284,-5310,13254,-5236 $DEVICE_ID=1003
MM673 VDD! 214 213 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12276 $Y=-3012  $PIN_XY=12306,-2940,12276,-3012,12246,-2940 $DEVICE_ID=1003
MM674 VDD! 182 181 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12276 $Y=-4160  $PIN_XY=12306,-4088,12276,-4160,12246,-4088 $DEVICE_ID=1003
MM675 VDD! 150 149 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12276 $Y=-5310  $PIN_XY=12306,-5236,12276,-5310,12246,-5236 $DEVICE_ID=1003
MM676 214 213 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11940 $Y=-3012  $PIN_XY=11970,-2940,11940,-3012,11910,-2940 $DEVICE_ID=1003
MM677 182 181 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11940 $Y=-4160  $PIN_XY=11970,-4088,11940,-4160,11910,-4088 $DEVICE_ID=1003
MM678 150 149 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11940 $Y=-5310  $PIN_XY=11970,-5236,11940,-5310,11910,-5236 $DEVICE_ID=1003
MM679 VDD! 212 211 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10932 $Y=-3012  $PIN_XY=10962,-2940,10932,-3012,10902,-2940 $DEVICE_ID=1003
MM680 VDD! 180 179 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10932 $Y=-4160  $PIN_XY=10962,-4088,10932,-4160,10902,-4088 $DEVICE_ID=1003
MM681 VDD! 148 147 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10932 $Y=-5310  $PIN_XY=10962,-5236,10932,-5310,10902,-5236 $DEVICE_ID=1003
MM682 212 211 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10596 $Y=-3012  $PIN_XY=10626,-2940,10596,-3012,10566,-2940 $DEVICE_ID=1003
MM683 180 179 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10596 $Y=-4160  $PIN_XY=10626,-4088,10596,-4160,10566,-4088 $DEVICE_ID=1003
MM684 148 147 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10596 $Y=-5310  $PIN_XY=10626,-5236,10596,-5310,10566,-5236 $DEVICE_ID=1003
MM685 VDD! 210 209 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9588 $Y=-3012  $PIN_XY=9618,-2940,9588,-3012,9558,-2940 $DEVICE_ID=1003
MM686 VDD! 178 177 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9588 $Y=-4160  $PIN_XY=9618,-4088,9588,-4160,9558,-4088 $DEVICE_ID=1003
MM687 VDD! 146 145 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9588 $Y=-5310  $PIN_XY=9618,-5236,9588,-5310,9558,-5236 $DEVICE_ID=1003
MM688 210 209 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9252 $Y=-3012  $PIN_XY=9282,-2940,9252,-3012,9222,-2940 $DEVICE_ID=1003
MM689 178 177 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9252 $Y=-4160  $PIN_XY=9282,-4088,9252,-4160,9222,-4088 $DEVICE_ID=1003
MM690 146 145 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9252 $Y=-5310  $PIN_XY=9282,-5236,9252,-5310,9222,-5236 $DEVICE_ID=1003
MM691 VDD! 208 207 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8244 $Y=-3012  $PIN_XY=8274,-2940,8244,-3012,8214,-2940 $DEVICE_ID=1003
MM692 VDD! 176 175 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8244 $Y=-4160  $PIN_XY=8274,-4088,8244,-4160,8214,-4088 $DEVICE_ID=1003
MM693 VDD! 144 143 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8244 $Y=-5310  $PIN_XY=8274,-5236,8244,-5310,8214,-5236 $DEVICE_ID=1003
MM694 208 207 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7908 $Y=-3012  $PIN_XY=7938,-2940,7908,-3012,7878,-2940 $DEVICE_ID=1003
MM695 176 175 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7908 $Y=-4160  $PIN_XY=7938,-4088,7908,-4160,7878,-4088 $DEVICE_ID=1003
MM696 144 143 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7908 $Y=-5310  $PIN_XY=7938,-5236,7908,-5310,7878,-5236 $DEVICE_ID=1003
MM697 VDD! 206 205 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6900 $Y=-3012  $PIN_XY=6930,-2940,6900,-3012,6870,-2940 $DEVICE_ID=1003
MM698 VDD! 174 173 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6900 $Y=-4160  $PIN_XY=6930,-4088,6900,-4160,6870,-4088 $DEVICE_ID=1003
MM699 VDD! 142 141 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6900 $Y=-5310  $PIN_XY=6930,-5236,6900,-5310,6870,-5236 $DEVICE_ID=1003
MM700 206 205 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6564 $Y=-3012  $PIN_XY=6594,-2940,6564,-3012,6534,-2940 $DEVICE_ID=1003
MM701 174 173 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6564 $Y=-4160  $PIN_XY=6594,-4088,6564,-4160,6534,-4088 $DEVICE_ID=1003
MM702 142 141 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6564 $Y=-5310  $PIN_XY=6594,-5236,6564,-5310,6534,-5236 $DEVICE_ID=1003
MM703 VDD! 204 203 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5556 $Y=-3012  $PIN_XY=5586,-2940,5556,-3012,5526,-2940 $DEVICE_ID=1003
MM704 VDD! 172 171 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5556 $Y=-4160  $PIN_XY=5586,-4088,5556,-4160,5526,-4088 $DEVICE_ID=1003
MM705 VDD! 140 139 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5556 $Y=-5310  $PIN_XY=5586,-5236,5556,-5310,5526,-5236 $DEVICE_ID=1003
MM706 204 203 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5220 $Y=-3012  $PIN_XY=5250,-2940,5220,-3012,5190,-2940 $DEVICE_ID=1003
MM707 172 171 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5220 $Y=-4160  $PIN_XY=5250,-4088,5220,-4160,5190,-4088 $DEVICE_ID=1003
MM708 140 139 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5220 $Y=-5310  $PIN_XY=5250,-5236,5220,-5310,5190,-5236 $DEVICE_ID=1003
MM709 VDD! 202 201 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4212 $Y=-3012  $PIN_XY=4242,-2940,4212,-3012,4182,-2940 $DEVICE_ID=1003
MM710 VDD! 170 169 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4212 $Y=-4160  $PIN_XY=4242,-4088,4212,-4160,4182,-4088 $DEVICE_ID=1003
MM711 VDD! 138 137 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4212 $Y=-5310  $PIN_XY=4242,-5236,4212,-5310,4182,-5236 $DEVICE_ID=1003
MM712 202 201 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3876 $Y=-3012  $PIN_XY=3906,-2940,3876,-3012,3846,-2940 $DEVICE_ID=1003
MM713 170 169 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3876 $Y=-4160  $PIN_XY=3906,-4088,3876,-4160,3846,-4088 $DEVICE_ID=1003
MM714 138 137 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3876 $Y=-5310  $PIN_XY=3906,-5236,3876,-5310,3846,-5236 $DEVICE_ID=1003
MM715 VDD! 200 199 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2868 $Y=-3012  $PIN_XY=2898,-2940,2868,-3012,2838,-2940 $DEVICE_ID=1003
MM716 VDD! 168 167 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2868 $Y=-4160  $PIN_XY=2898,-4088,2868,-4160,2838,-4088 $DEVICE_ID=1003
MM717 VDD! 136 135 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2868 $Y=-5310  $PIN_XY=2898,-5236,2868,-5310,2838,-5236 $DEVICE_ID=1003
MM718 200 199 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2532 $Y=-3012  $PIN_XY=2562,-2940,2532,-3012,2502,-2940 $DEVICE_ID=1003
MM719 168 167 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2532 $Y=-4160  $PIN_XY=2562,-4088,2532,-4160,2502,-4088 $DEVICE_ID=1003
MM720 136 135 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2532 $Y=-5310  $PIN_XY=2562,-5236,2532,-5310,2502,-5236 $DEVICE_ID=1003
MM721 VDD! 198 197 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1524 $Y=-3012  $PIN_XY=1554,-2940,1524,-3012,1494,-2940 $DEVICE_ID=1003
MM722 VDD! 166 165 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1524 $Y=-4160  $PIN_XY=1554,-4088,1524,-4160,1494,-4088 $DEVICE_ID=1003
MM723 VDD! 134 133 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1524 $Y=-5310  $PIN_XY=1554,-5236,1524,-5310,1494,-5236 $DEVICE_ID=1003
MM724 198 197 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1188 $Y=-3012  $PIN_XY=1218,-2940,1188,-3012,1158,-2940 $DEVICE_ID=1003
MM725 166 165 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1188 $Y=-4160  $PIN_XY=1218,-4088,1188,-4160,1158,-4088 $DEVICE_ID=1003
MM726 134 133 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1188 $Y=-5310  $PIN_XY=1218,-5236,1188,-5310,1158,-5236 $DEVICE_ID=1003
MM727 VDD! 196 195 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=180 $Y=-3012  $PIN_XY=210,-2940,180,-3012,150,-2940 $DEVICE_ID=1003
MM728 VDD! 164 163 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=180 $Y=-4160  $PIN_XY=210,-4088,180,-4160,150,-4088 $DEVICE_ID=1003
MM729 VDD! 132 131 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=180 $Y=-5310  $PIN_XY=210,-5236,180,-5310,150,-5236 $DEVICE_ID=1003
MM730 196 195 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=-156 $Y=-3012  $PIN_XY=-126,-2940,-156,-3012,-186,-2940 $DEVICE_ID=1003
MM731 164 163 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=-156 $Y=-4160  $PIN_XY=-126,-4088,-156,-4160,-186,-4088 $DEVICE_ID=1003
MM732 132 131 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=-156 $Y=-5310  $PIN_XY=-126,-5236,-156,-5310,-186,-5236 $DEVICE_ID=1003
MM733 VDD! 130 129 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20340 $Y=-6457  $PIN_XY=20370,-6382,20340,-6457,20310,-6382 $DEVICE_ID=1003
MM734 VDD! 98 97 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20340 $Y=-7581  $PIN_XY=20370,-7530,20340,-7581,20310,-7530 $DEVICE_ID=1003
MM735 130 129 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20004 $Y=-6457  $PIN_XY=20034,-6382,20004,-6457,19974,-6382 $DEVICE_ID=1003
MM736 98 97 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=20004 $Y=-7581  $PIN_XY=20034,-7530,20004,-7581,19974,-7530 $DEVICE_ID=1003
MM737 VDD! 128 127 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18996 $Y=-6457  $PIN_XY=19026,-6382,18996,-6457,18966,-6382 $DEVICE_ID=1003
MM738 VDD! 96 95 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18996 $Y=-7596  $PIN_XY=19026,-7530,18996,-7596,18966,-7530 $DEVICE_ID=1003
MM739 128 127 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18660 $Y=-6457  $PIN_XY=18690,-6382,18660,-6457,18630,-6382 $DEVICE_ID=1003
MM740 96 95 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=18660 $Y=-7581  $PIN_XY=18690,-7530,18660,-7581,18630,-7530 $DEVICE_ID=1003
MM741 VDD! 126 125 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17652 $Y=-6457  $PIN_XY=17682,-6382,17652,-6457,17622,-6382 $DEVICE_ID=1003
MM742 VDD! 94 93 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17652 $Y=-7581  $PIN_XY=17682,-7530,17652,-7581,17622,-7530 $DEVICE_ID=1003
MM743 126 125 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17316 $Y=-6457  $PIN_XY=17346,-6382,17316,-6457,17286,-6382 $DEVICE_ID=1003
MM744 94 93 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=17316 $Y=-7581  $PIN_XY=17346,-7530,17316,-7581,17286,-7530 $DEVICE_ID=1003
MM745 VDD! 124 123 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16308 $Y=-6457  $PIN_XY=16338,-6382,16308,-6457,16278,-6382 $DEVICE_ID=1003
MM746 VDD! 92 91 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=16308 $Y=-7581  $PIN_XY=16338,-7530,16308,-7581,16278,-7530 $DEVICE_ID=1003
MM747 124 123 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15972 $Y=-6457  $PIN_XY=16002,-6382,15972,-6457,15942,-6382 $DEVICE_ID=1003
MM748 92 91 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=15972 $Y=-7581  $PIN_XY=16002,-7530,15972,-7581,15942,-7530 $DEVICE_ID=1003
MM749 VDD! 122 121 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14964 $Y=-6457  $PIN_XY=14994,-6382,14964,-6457,14934,-6382 $DEVICE_ID=1003
MM750 VDD! 90 89 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14964 $Y=-7581  $PIN_XY=14994,-7530,14964,-7581,14934,-7530 $DEVICE_ID=1003
MM751 122 121 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14628 $Y=-6457  $PIN_XY=14658,-6382,14628,-6457,14598,-6382 $DEVICE_ID=1003
MM752 90 89 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=14628 $Y=-7581  $PIN_XY=14658,-7530,14628,-7581,14598,-7530 $DEVICE_ID=1003
MM753 VDD! 120 119 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13620 $Y=-6457  $PIN_XY=13650,-6382,13620,-6457,13590,-6382 $DEVICE_ID=1003
MM754 VDD! 88 87 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13620 $Y=-7596  $PIN_XY=13650,-7530,13620,-7596,13590,-7530 $DEVICE_ID=1003
MM755 120 119 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13284 $Y=-6457  $PIN_XY=13314,-6382,13284,-6457,13254,-6382 $DEVICE_ID=1003
MM756 88 87 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=13284 $Y=-7581  $PIN_XY=13314,-7530,13284,-7581,13254,-7530 $DEVICE_ID=1003
MM757 VDD! 118 117 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12276 $Y=-6457  $PIN_XY=12306,-6382,12276,-6457,12246,-6382 $DEVICE_ID=1003
MM758 VDD! 86 85 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=12276 $Y=-7581  $PIN_XY=12306,-7530,12276,-7581,12246,-7530 $DEVICE_ID=1003
MM759 118 117 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11940 $Y=-6457  $PIN_XY=11970,-6382,11940,-6457,11910,-6382 $DEVICE_ID=1003
MM760 86 85 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=11940 $Y=-7581  $PIN_XY=11970,-7530,11940,-7581,11910,-7530 $DEVICE_ID=1003
MM761 VDD! 116 115 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10932 $Y=-6457  $PIN_XY=10962,-6382,10932,-6457,10902,-6382 $DEVICE_ID=1003
MM762 VDD! 84 83 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10932 $Y=-7581  $PIN_XY=10962,-7530,10932,-7581,10902,-7530 $DEVICE_ID=1003
MM763 116 115 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10596 $Y=-6457  $PIN_XY=10626,-6382,10596,-6457,10566,-6382 $DEVICE_ID=1003
MM764 84 83 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=10596 $Y=-7581  $PIN_XY=10626,-7530,10596,-7581,10566,-7530 $DEVICE_ID=1003
MM765 VDD! 114 113 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9588 $Y=-6457  $PIN_XY=9618,-6382,9588,-6457,9558,-6382 $DEVICE_ID=1003
MM766 VDD! 82 81 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9588 $Y=-7581  $PIN_XY=9618,-7530,9588,-7581,9558,-7530 $DEVICE_ID=1003
MM767 114 113 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9252 $Y=-6457  $PIN_XY=9282,-6382,9252,-6457,9222,-6382 $DEVICE_ID=1003
MM768 82 81 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=9252 $Y=-7581  $PIN_XY=9282,-7530,9252,-7581,9222,-7530 $DEVICE_ID=1003
MM769 VDD! 112 111 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8244 $Y=-6457  $PIN_XY=8274,-6382,8244,-6457,8214,-6382 $DEVICE_ID=1003
MM770 VDD! 80 79 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=8244 $Y=-7581  $PIN_XY=8274,-7530,8244,-7581,8214,-7530 $DEVICE_ID=1003
MM771 112 111 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7908 $Y=-6457  $PIN_XY=7938,-6382,7908,-6457,7878,-6382 $DEVICE_ID=1003
MM772 80 79 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=7908 $Y=-7581  $PIN_XY=7938,-7530,7908,-7581,7878,-7530 $DEVICE_ID=1003
MM773 VDD! 110 109 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6900 $Y=-6457  $PIN_XY=6930,-6382,6900,-6457,6870,-6382 $DEVICE_ID=1003
MM774 VDD! 78 77 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6900 $Y=-7581  $PIN_XY=6930,-7530,6900,-7581,6870,-7530 $DEVICE_ID=1003
MM775 110 109 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6564 $Y=-6457  $PIN_XY=6594,-6382,6564,-6457,6534,-6382 $DEVICE_ID=1003
MM776 78 77 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=6564 $Y=-7581  $PIN_XY=6594,-7530,6564,-7581,6534,-7530 $DEVICE_ID=1003
MM777 VDD! 108 107 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5556 $Y=-6457  $PIN_XY=5586,-6382,5556,-6457,5526,-6382 $DEVICE_ID=1003
MM778 VDD! 76 75 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5556 $Y=-7581  $PIN_XY=5586,-7530,5556,-7581,5526,-7530 $DEVICE_ID=1003
MM779 108 107 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5220 $Y=-6457  $PIN_XY=5250,-6382,5220,-6457,5190,-6382 $DEVICE_ID=1003
MM780 76 75 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=5220 $Y=-7581  $PIN_XY=5250,-7530,5220,-7581,5190,-7530 $DEVICE_ID=1003
MM781 VDD! 106 105 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4212 $Y=-6457  $PIN_XY=4242,-6382,4212,-6457,4182,-6382 $DEVICE_ID=1003
MM782 VDD! 74 73 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=4212 $Y=-7581  $PIN_XY=4242,-7530,4212,-7581,4182,-7530 $DEVICE_ID=1003
MM783 106 105 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3876 $Y=-6457  $PIN_XY=3906,-6382,3876,-6457,3846,-6382 $DEVICE_ID=1003
MM784 74 73 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=3876 $Y=-7581  $PIN_XY=3906,-7530,3876,-7581,3846,-7530 $DEVICE_ID=1003
MM785 VDD! 104 103 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2868 $Y=-6457  $PIN_XY=2898,-6382,2868,-6457,2838,-6382 $DEVICE_ID=1003
MM786 VDD! 72 71 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2868 $Y=-7581  $PIN_XY=2898,-7530,2868,-7581,2838,-7530 $DEVICE_ID=1003
MM787 104 103 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2532 $Y=-6457  $PIN_XY=2562,-6382,2532,-6457,2502,-6382 $DEVICE_ID=1003
MM788 72 71 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=2532 $Y=-7581  $PIN_XY=2562,-7530,2532,-7581,2502,-7530 $DEVICE_ID=1003
MM789 VDD! 102 101 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1524 $Y=-6457  $PIN_XY=1554,-6382,1524,-6457,1494,-6382 $DEVICE_ID=1003
MM790 VDD! 70 69 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1524 $Y=-7581  $PIN_XY=1554,-7530,1524,-7581,1494,-7530 $DEVICE_ID=1003
MM791 102 101 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1188 $Y=-6457  $PIN_XY=1218,-6382,1188,-6457,1158,-6382 $DEVICE_ID=1003
MM792 70 69 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=1188 $Y=-7581  $PIN_XY=1218,-7530,1188,-7581,1158,-7530 $DEVICE_ID=1003
MM793 VDD! 100 99 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=180 $Y=-6457  $PIN_XY=210,-6382,180,-6457,150,-6382 $DEVICE_ID=1003
MM794 VDD! 68 67 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=180 $Y=-7581  $PIN_XY=210,-7530,180,-7581,150,-7530 $DEVICE_ID=1003
MM795 100 99 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=-156 $Y=-6457  $PIN_XY=-126,-6382,-156,-6457,-186,-6382 $DEVICE_ID=1003
MM796 68 67 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=-156 $Y=-7581  $PIN_XY=-126,-7530,-156,-7581,-186,-7530 $DEVICE_ID=1003
MM797 333 332 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=23534 $Y=-20675  $PIN_XY=23564,-20698,23534,-20675,23504,-20698 $DEVICE_ID=1003
MM798 332 CLK VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=23198 $Y=-20678  $PIN_XY=23228,-20698,23198,-20678,23168,-20698 $DEVICE_ID=1003
MM799 331 CLK 1535 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=22862 $Y=-20696  $PIN_XY=22892,-20698,22862,-20696,22832,-20698 $DEVICE_ID=1003
MM800 1535 2 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=22694 $Y=-20696  $PIN_XY=22724,-20698,22694,-20696,22664,-20698 $DEVICE_ID=1003
MM801 Q<0> 334 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=24374 $Y=-20862  $PIN_XY=(24404,-20698,24404,-20868),24374,-20862,(24344,-20698,24344,-20868) $DEVICE_ID=1003
MM802 Q<1> 330 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=24374 $Y=-22750  $PIN_XY=(24404,-22586,24404,-22756),24374,-22750,(24344,-22586,24344,-22756) $DEVICE_ID=1003
MM803 334 333 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=24038 $Y=-20863  $PIN_XY=(24068,-20698,24068,-20868),24038,-20863,(24008,-20698,24008,-20868) $DEVICE_ID=1003
MM804 330 329 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=24038 $Y=-22751  $PIN_XY=(24068,-22586,24068,-22756),24038,-22751,(24008,-22586,24008,-22756) $DEVICE_ID=1003
MM805 329 328 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=23534 $Y=-22563  $PIN_XY=23564,-22586,23534,-22563,23504,-22586 $DEVICE_ID=1003
MM806 337 336 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=23534 $Y=-24451  $PIN_XY=23564,-24474,23534,-24451,23504,-24474 $DEVICE_ID=1003
MM807 328 CLK VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=23198 $Y=-22566  $PIN_XY=23228,-22586,23198,-22566,23168,-22586 $DEVICE_ID=1003
MM808 336 CLK VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=23198 $Y=-24454  $PIN_XY=23228,-24474,23198,-24454,23168,-24474 $DEVICE_ID=1003
MM809 327 CLK 1534 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=22862 $Y=-22584  $PIN_XY=22892,-22586,22862,-22584,22832,-22586 $DEVICE_ID=1003
MM810 1534 4 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=22694 $Y=-22584  $PIN_XY=22724,-22586,22694,-22584,22664,-22586 $DEVICE_ID=1003
MM811 Q<2> 338 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=24374 $Y=-24638  $PIN_XY=(24404,-24474,24404,-24644),24374,-24638,(24344,-24474,24344,-24644) $DEVICE_ID=1003
MM812 Q<3> 326 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=24374 $Y=-26526  $PIN_XY=(24404,-26362,24404,-26532),24374,-26526,(24344,-26362,24344,-26532) $DEVICE_ID=1003
MM813 338 337 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=24038 $Y=-24639  $PIN_XY=(24068,-24474,24068,-24644),24038,-24639,(24008,-24474,24008,-24644) $DEVICE_ID=1003
MM814 326 325 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=4 ADEO=5.67e-16 ASEO=5.67e-16 PDEO=1.17e-07
+	 PSEO=1.17e-07 $X=24038 $Y=-26527  $PIN_XY=(24068,-26362,24068,-26532),24038,-26527,(24008,-26362,24008,-26532) $DEVICE_ID=1003
MM815 325 324 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=23534 $Y=-26339  $PIN_XY=23564,-26362,23534,-26339,23504,-26362 $DEVICE_ID=1003
MM816 324 CLK VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=2.835e-16 PDEO=5.85e-08
+	 PSEO=5.85e-08 $X=23198 $Y=-26342  $PIN_XY=23228,-26362,23198,-26342,23168,-26362 $DEVICE_ID=1003
MM817 335 CLK 1536 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=22862 $Y=-24472  $PIN_XY=22892,-24474,22862,-24472,22832,-24474 $DEVICE_ID=1003
MM818 323 CLK 1533 pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=2.835e-16 ASEO=5.67e-16 PDEO=5.85e-08
+	 PSEO=1.17e-07 $X=22862 $Y=-26360  $PIN_XY=22892,-26362,22862,-26360,22832,-26362 $DEVICE_ID=1003
MM819 1536 8 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=22694 $Y=-24472  $PIN_XY=22724,-24474,22694,-24472,22664,-24474 $DEVICE_ID=1003
MM820 1533 6 VDD! pmos  W=2.1e-08 L=1.5e-08 NFIN=2 ADEO=5.67e-16 ASEO=2.835e-16 PDEO=1.17e-07
+	 PSEO=5.85e-08 $X=22694 $Y=-26360  $PIN_XY=22724,-26362,22694,-26360,22664,-26362 $DEVICE_ID=1003
XX880FE34C1 12 13 CLK 15 16 CLK VDD! GND! VDD! GND! 1521 
+	VDD! VDD! VCELLR2 $T=-2654 3310 0 0 $X=-548 $Y=4658
XX880FE34C2 17 18 CLK 19 20 CLK VDD! GND! VDD! GND! 1521 
+	VDD! VDD! VCELLR2 $T=-638 3310 0 0 $X=1468 $Y=4658
XX880FE34C3 21 22 CLK 23 24 CLK VDD! GND! VDD! GND! 1521 
+	VDD! VDD! VCELLR2 $T=2722 3310 0 0 $X=4827 $Y=4658
XX880FE34C4 25 26 CLK 27 28 CLK VDD! GND! VDD! GND! 1521 
+	VDD! VDD! VCELLR2 $T=4738 3310 0 0 $X=6844 $Y=4658
XX880FE34C5 29 30 CLK 31 32 CLK VDD! GND! VDD! GND! 1521 
+	VDD! VDD! VCELLR2 $T=8098 3310 0 0 $X=10204 $Y=4658
XX880FE34C6 33 34 CLK 35 36 CLK VDD! GND! VDD! GND! 1521 
+	VDD! VDD! VCELLR2 $T=10114 3310 0 0 $X=12220 $Y=4658
XX880FE34C7 37 38 CLK 39 40 CLK VDD! GND! VDD! GND! 1521 
+	VDD! VDD! VCELLR2 $T=13474 3310 0 0 $X=15580 $Y=4658
XX880FE34C8 41 42 CLK 43 44 CLK VDD! GND! VDD! GND! 1521 
+	VDD! VDD! VCELLR2 $T=15490 3310 0 0 $X=17596 $Y=4658
XX880FE34C9 2 3 D<0> WENB GND! VDD! 1522 VDD! VDD! VDD! GND! Write_Driver $T=598 -30806 0 0 $X=20 $Y=-30782
XX880FE34C10 4 5 D<1> WENB GND! VDD! 1522 VDD! VDD! 1531 1537 Write_Driver $T=6312 -30806 0 0 $X=5734 $Y=-30782
XX880FE34C11 6 7 D<3> WENB GND! VDD! 1522 VDD! VDD! VDD! GND! Write_Driver $T=17742 -30806 0 0 $X=17164 $Y=-30782
XX880FE34C12 8 9 D<2> WENB GND! VDD! 1522 VDD! VDD! 1532 1538 Write_Driver $T=12028 -30806 0 0 $X=11450 $Y=-30782
XX880FE34C13 A<3> VDD! A<4> GND! A<2> 60 59 58 57 56 55 
+	54 53 rowdecoder $T=-17680 -8206 0 0 $X=-17534 $Y=-8071
XX880FE34C14 A<0> A<1> 16 18 20 12 15 17 19 22 24 
+	26 28 21 23 25 27 30 32 34 36 29 
+	31 33 35 38 40 42 44 37 39 41 43 
+	2 13 4 8 6 3 5 9 7 VDD! GND! 
+	VDD! column_decoder_new $T=7500 -16254 0 0 $X=564 $Y=-19206
XX880FE34C15 53 53 53 53 53 53 53 53 67 68 69 
+	70 71 72 73 74 75 76 77 78 79 80 
+	81 82 339 340 341 342 343 344 345 346 347 
+	348 349 350 351 352 353 354 GND! VDD! GND! VDD! 
+	GND! VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! VDD! 
+	GND! 12 13 15 16 17 18 19 20 21 22 
+	23 24 25 26 27 28 1524 VDD! VCELLR4 $T=-156 -7700 0 0 $X=-714 $Y=-8109
XX880FE34C16 53 53 53 53 53 53 53 53 83 84 85 
+	86 87 88 89 90 91 92 93 94 95 96 
+	97 98 355 356 357 358 359 360 361 362 363 
+	364 365 366 367 368 369 370 GND! VDD! GND! VDD! 
+	GND! VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! VDD! 
+	GND! 29 30 31 32 33 34 35 36 37 38 
+	39 40 41 42 43 44 1524 VDD! VCELLR4 $T=10596 -7700 0 0 $X=10038 $Y=-8109
XX880FE34C17 54 54 54 54 54 54 54 54 99 100 101 
+	102 103 104 105 106 107 108 109 110 111 112 
+	113 114 371 372 373 374 375 376 377 378 379 
+	380 381 382 383 384 385 386 GND! VDD! GND! VDD! 
+	GND! VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! VDD! 
+	GND! 12 13 15 16 17 18 19 20 21 22 
+	23 24 25 26 27 28 1525 VDD! VCELLR4 $T=-156 -6552 0 0 $X=-714 $Y=-6962
XX880FE34C18 54 54 54 54 54 54 54 54 115 116 117 
+	118 119 120 121 122 123 124 125 126 127 128 
+	129 130 387 388 389 390 391 392 393 394 395 
+	396 397 398 399 400 401 402 GND! VDD! GND! VDD! 
+	GND! VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! VDD! 
+	GND! 29 30 31 32 33 34 35 36 37 38 
+	39 40 41 42 43 44 1525 VDD! VCELLR4 $T=10596 -6552 0 0 $X=10038 $Y=-6962
XX880FE34C19 55 55 55 55 55 55 55 55 131 132 133 
+	134 135 136 137 138 139 140 141 142 143 144 
+	145 146 403 404 405 406 407 408 409 410 411 
+	412 413 414 415 416 417 418 GND! VDD! GND! VDD! 
+	GND! VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! VDD! 
+	GND! 12 13 15 16 17 18 19 20 21 22 
+	23 24 25 26 27 28 1526 VDD! VCELLR4 $T=-156 -5406 0 0 $X=-714 $Y=-5816
XX880FE34C20 55 55 55 55 55 55 55 55 147 148 149 
+	150 151 152 153 154 155 156 157 158 159 160 
+	161 162 419 420 421 422 423 424 425 426 427 
+	428 429 430 431 432 433 434 GND! VDD! GND! VDD! 
+	GND! VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! VDD! 
+	GND! 29 30 31 32 33 34 35 36 37 38 
+	39 40 41 42 43 44 1526 VDD! VCELLR4 $T=10596 -5406 0 0 $X=10038 $Y=-5816
XX880FE34C21 56 56 56 56 56 56 56 56 163 164 165 
+	166 167 168 169 170 171 172 173 174 175 176 
+	177 178 435 436 437 438 439 440 441 442 443 
+	444 445 446 447 448 449 450 GND! VDD! GND! VDD! 
+	GND! VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! VDD! 
+	GND! 12 13 15 16 17 18 19 20 21 22 
+	23 24 25 26 27 28 1527 VDD! VCELLR4 $T=-156 -4258 0 0 $X=-714 $Y=-4668
XX880FE34C22 56 56 56 56 56 56 56 56 179 180 181 
+	182 183 184 185 186 187 188 189 190 191 192 
+	193 194 451 452 453 454 455 456 457 458 459 
+	460 461 462 463 464 465 466 GND! VDD! GND! VDD! 
+	GND! VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! VDD! 
+	GND! 29 30 31 32 33 34 35 36 37 38 
+	39 40 41 42 43 44 1527 VDD! VCELLR4 $T=10596 -4258 0 0 $X=10038 $Y=-4668
XX880FE34C23 57 57 57 57 57 57 57 57 195 196 197 
+	198 199 200 201 202 203 204 205 206 207 208 
+	209 210 467 468 469 470 471 472 473 474 475 
+	476 477 478 479 480 481 482 GND! VDD! GND! VDD! 
+	GND! VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! VDD! 
+	GND! 12 13 15 16 17 18 19 20 21 22 
+	23 24 25 26 27 28 1528 VDD! VCELLR4 $T=-156 -3110 0 0 $X=-714 $Y=-3520
XX880FE34C24 57 57 57 57 57 57 57 57 211 212 213 
+	214 215 216 217 218 219 220 221 222 223 224 
+	225 226 483 484 485 486 487 488 489 490 491 
+	492 493 494 495 496 497 498 GND! VDD! GND! VDD! 
+	GND! VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! VDD! 
+	GND! 29 30 31 32 33 34 35 36 37 38 
+	39 40 41 42 43 44 1528 VDD! VCELLR4 $T=10596 -3110 0 0 $X=10038 $Y=-3520
XX880FE34C25 58 58 58 58 58 58 58 58 227 228 229 
+	230 231 232 233 234 235 236 237 238 239 240 
+	241 242 499 500 501 502 503 504 505 506 507 
+	508 509 510 511 512 513 514 GND! VDD! GND! VDD! 
+	GND! VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! VDD! 
+	GND! 12 13 15 16 17 18 19 20 21 22 
+	23 24 25 26 27 28 1529 VDD! VCELLR4 $T=-156 -1962 0 0 $X=-714 $Y=-2372
XX880FE34C26 58 58 58 58 58 58 58 58 243 244 245 
+	246 247 248 249 250 251 252 253 254 255 256 
+	257 258 515 516 517 518 519 520 521 522 523 
+	524 525 526 527 528 529 530 GND! VDD! GND! VDD! 
+	GND! VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! VDD! 
+	GND! 29 30 31 32 33 34 35 36 37 38 
+	39 40 41 42 43 44 1529 VDD! VCELLR4 $T=10596 -1962 0 0 $X=10038 $Y=-2372
XX880FE34C27 59 59 59 59 59 59 59 59 259 260 261 
+	262 263 264 265 266 267 268 269 270 271 272 
+	273 274 531 532 533 534 535 536 537 538 539 
+	540 541 542 543 544 545 546 GND! VDD! GND! VDD! 
+	GND! VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! VDD! 
+	GND! 12 13 15 16 17 18 19 20 21 22 
+	23 24 25 26 27 28 1530 VDD! VCELLR4 $T=-156 -816 0 0 $X=-714 $Y=-1226
XX880FE34C28 59 59 59 59 59 59 59 59 275 276 277 
+	278 279 280 281 282 283 284 285 286 287 288 
+	289 290 547 548 549 550 551 552 553 554 555 
+	556 557 558 559 560 561 562 GND! VDD! GND! VDD! 
+	GND! VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! VDD! 
+	GND! 29 30 31 32 33 34 35 36 37 38 
+	39 40 41 42 43 44 1530 VDD! VCELLR4 $T=10596 -816 0 0 $X=10038 $Y=-1226
XX880FE34C29 60 60 60 60 60 60 60 60 291 292 293 
+	294 295 296 297 298 299 300 301 302 303 304 
+	305 306 563 564 565 566 567 568 569 570 571 
+	572 573 574 575 576 577 578 GND! VDD! GND! VDD! 
+	GND! VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! VDD! 
+	GND! 12 13 15 16 17 18 19 20 21 22 
+	23 24 25 26 27 28 1523 VDD! VCELLR4 $T=-156 332 0 0 $X=-714 $Y=-78
XX880FE34C30 60 60 60 60 60 60 60 60 307 308 309 
+	310 311 312 313 314 315 316 317 318 319 320 
+	321 322 579 580 581 582 583 584 585 586 587 
+	588 589 590 591 592 593 594 GND! VDD! GND! VDD! 
+	GND! VDD! GND! VDD! GND! VDD! VDD! GND! VDD! GND! VDD! 
+	GND! 29 30 31 32 33 34 35 36 37 38 
+	39 40 41 42 43 44 1523 VDD! VCELLR4 $T=10596 332 0 0 $X=10038 $Y=-78
XX880FE34C31 6 323 CLK 324 Q<3> 325 326 GND! VDD! 1533 1539 
+	1540 VDD! VDD! tspc_flip_flop $T=20916 -27794 0 0 $X=22472 $Y=-27090
XX880FE34C32 4 327 CLK 328 Q<1> 329 330 GND! VDD! 1534 1541 
+	1542 VDD! VDD! tspc_flip_flop $T=20916 -24018 0 0 $X=22472 $Y=-23314
XX880FE34C33 2 331 CLK 332 Q<0> 333 334 GND! VDD! 1535 1543 
+	1544 VDD! VDD! tspc_flip_flop $T=20916 -22130 0 0 $X=22472 $Y=-21426
XX880FE34C34 8 335 CLK 336 Q<2> 337 338 GND! VDD! 1536 1545 
+	1546 VDD! VDD! tspc_flip_flop $T=20916 -25906 0 0 $X=22472 $Y=-25202
.ends bit_cell_array
